XlxV64EB    fa00    2700o���i���y���O㓕�Dh0��숤?L8�A��`a���ʸ+"��/�o� �D�z=��W��UW'DjK�V�\	�'�~'$�<M�{I��Ab0%U�+�����;�S{�ɘ��hc��1��Lu=�j}�`�FmhFy�ݠ��g�QY�T��P�k%�A�H�_AmT���"�<}|��᎝s3�45�B�"�>�;�.۶!��ٸ-q)R6CW�Ǻ!e2�.�1p�#�q=3����[��5Rs]bhx^��XlX�;��-U���i)�����Ow�G�/���̄����~�%h|��*0��8Im���xMp�\[K.������
�[�EҘ�P�.��4�����T��WͿHx���ѼK�\� �/�B\�[�ݨ�t��f��ܱ](?� ��4>g�%�zb�G����~'�D�Z�k ��5�Y��-ǡWY�����fK��V=QZ�4�=�5���T&������#�R�A�5:���}e��1"W	���V ���O��,����"�0o��!Mxq���7.�I�D�^��4�,�$�Q ;\�.-�4��Y��ږ��xM���z���>���v�4jI������<��S���r���Ѧ_aI��L��wN������' w��DB�n�ϱ{Y��s��Js�Too�<즤�O"L'z�����q��e&[=' "�,v�t��#$s!ѹ�|"���-�}�2N���� ��C�z*G/c����I��M�E��n�`S�I���eJB6
{�b~p'T��(='�n2��I������ݵ�{��������,���Occp���A�
�n�R2����0lEo�I��F�Y�t3�u�J@fe�P���)�!(�l"���\7A�繅Y��S{�t����j�3��8�D�d���^{Бk���p�A�
����Y@ݡ]��Z;C�.:x����EQ(��G,<VzC�3�v;gu�T�#ip��˪x#����!�?q��c�shq�����ؤ�鏶}��F�$��=:�:$�� �����{����<Ђ�6]�����É0������Z��bˀh|�P����W�Wi��AZ]���;s��!�6P�|9nR%ƍ�J1Ϣ+�V�3C\����&�D����x����P�q@�]��Ƹ�8�`��ܞ7^�)t7p4�)�,���4Dd���CG��_`k����o-l]��i����Tm���tϟT�v����E}��J%�+:/U��~�N��>�;�i3���<���h���1Ұ��1(��1����%��z�U�]��/��rZ��_^O9G��.
X	�P��(���axݔ�9ka�w0��{�$p9�ߪr�j��w����[$~������x8���)HA|��nS5�}�+g����F2l6:
���YbL6!Epi�Ɩ<mŲ��n6�֭�gǉCě�=^#��� UrV�H��7��Z�WĆ�h~�9	c�cq<(�X��Н*��M�H��Y'~I�1�<;�\�Y�3�[��7��
C�q̂�o#q��p��^+ȭ��
�zg�n�f��s�:���K�@6�~��l@�Ywu��	/�Ys�6XW�w�LB��Cax�������fף�^`}��i�-F����],�����͜P,�WCU�["ZCڈ�euS(C�m�������j�ɤ(��@(��ǻ��x�/���nFt���$�c2��mno�H��U��`�U��E5��5��\J|��,��i�-Q.�l����_T�C��Lm�RA���u|������G�_��+Q�͠���Z�mm���\J]�{�X꺋m~�e�w)NĶ������"��/�n�;&��+���uG#G.��Qċ ��}٨��;�8hE��\c���1B���2V8�ža����$�5��Z��&Q�u�H����I)"��v�m������u%�����N�6��q��@�F���`�s�:�[�JTdg�#�I��U�J�ك"��xNa�����Pv��)z~aZ ���c��xOk�O'~p=���+���>�M:�_H�ƒ�9	�+��b��n0�	�G J�Y��6���Sa�W��E���s2�ݢ�p��At'��D��wA<��`1�fU!���P���G�c��V)?-��u��w��s������j�O�Z�Fmq��!���xd����K����Ui�+6>vC��[s �|����j�3���f�/�Q�,Uf�63�e�W ���'�[��lG�?��V�܀V�	(�R���R�T��*sj̱O�he��oq�}5�$�f��9��}<\��zp����`IZ�j�E*U���'���T�T[/V9�Jc��%!�t�Ga�.(S}�B���C�.����	sP'�'���q���o��o��x�!��R��C�~��E�8l�zUܼ�4���09�G�S�2tQ(��PO��ѭ�Y��)_Q�����μ��)�r�:�X�,ٹ����{�MC>�TA�#�������P��KUE�=\A�����<��P�R��z�5��[�9�Ds�v"$J�����Q��.\��k�J�7��#�����+�?���WI2Zl2sax����-"�Sܴ�*]��c�#�}7�D���R�R��._dO�pG�,���g�N[W���~���cF�wGF+ݴ� �����AL��`��,hL��bʖ0��:��7����od_�ne��/�b.�Bk��y�<N�E%='t!�Ty"�;	�����E��
�O!�7�u�[\��6`4!B�=����2��g��1�.�,��WՖ�8[3\�MW�F�����̈́�ċ��z`N�yI��L�t��J�V*��rF�\N�^xӧQ�!˨TǷB$�����,��Ъ������}g��V�wS����-�f�L��`�T)yqf�  �I.��xΝ8*Yf���?�@��I���1�;�i�D��}�`mM��-N�_b`�V
�pStN^�����Wu��>s���6�1e�|�#9p��CeX�/�:�K���7�.-=����ц>"{�f6s5���
��i����x�Kڱ1d��Kz87�[*_@��m�xH59|s�TCM�q��/���z��QExAw],[�Mcj���{T�d��/���+(5Ք��S;�4�t�/m�5���:�G٪=���?�-����J�" �p�-وT#=���q�;�?'{�]��oz@�+e�8�%�u��MAs՗���ޑ���^JGy�|.�x�9�M�u�l%bm����iw�G���}9��
�H.,��[���zy �c�+v�&>C
�(�����0@,�xVa�O1;0t��Zy7�K�-�\bF'qqZ꬙l�A��T7��~�}�lG(�nX�$��ஐv�_A��\\��=��iW��<J��f�
ł7��5�7Ӂ�/���h���`�T��7 ��Y�(n��No��������I�i�rx墳��F���γY�����s|�W�e<�n#\e5�N�18'�}�pi�G�l#'�֢��+��u� �o�hlB�|w�V�!��z:�gs�-~�2�O���\�zU�j��g�{An�e�U�|����IU���TP��i�|���%�Ki E��97�M�]�&U��:�OE�y�rmg��$,��9& �3g��됱gr8 "�qZ1M��3��S�>�
r�f͉m��ѝN��~�C�vB����t�
w0�1�)���j;Ƚ����8�j�f�P\5��0��D5A'�rU{|~
Z�?X�b�m��4&E�d ��.sm�I��o��U�y��?�M�v�i��Zc��*�c�]��0�j�C{��\���L�G�؍q#���uu�HG�3��pS�9ٻd�"~3�̡b���FP+����'J���daM7���<�>�سBψ"6�k$Sg��B˧���t�n�>�O.���l��}��u�D�v$�ܿ/��;�Z+����s�R:N̵���#�~v�8>�ݢ�b������BfH�Rݐ�5�����Ɇ�ʿ	g{�(Zr�s�Rm�8/�ߧ��(|�V@W�D&�� �cs��=��FP�?�6� �5qJL���Ǉ9�|�!�u�`i�
�s�P&A,N�N�>��Z:�t���F�5�CZ��, ��`qf ɥ�8  �ʗ&7f�"V�U����ӧ��F�^�m�n�;Ҵj�B�Z�T��P}��X�C~��Xh|\OyL��G�}�jx{By�C�`��j/��%|��4�pE�r��^�ޕ���!�Mt�R���ڐ�²M ����0��7��g�����;�
�"�lM�b�w�џ�J�ޅj��1B%�����6��Iz�v�����o���z���!p�"�:lq��?��������9�w9`aͰ�z΍���r��I!x�89@��p��f�o��K�ޞ�h/8*��>�R�r[��_���1ƒ���S���ŽV����v�!-���_�����=Z+�R����%l��1l��oμ0M;�3�8t[ƠEH3Sw�>�Ι��K����p�^+4�;Y��h��D��rK�h�a�!������'Z-����%��ȢN]�ы�8N80��5�k!A�{��%���"�E�O�P�[?��l��-h��ؖG;�@M$<Zr�Sx�*�(�&_�7��:��Cu����үL��1U2� �-�ɱ,���Z%�UD�j&{�n���s%]Ĥ��7��M3�>x����^�A����^�gָ?���"�铘|��>z���/�$|����\Iܜ䙊ȿB:��{��tBs����Y�w�R��U�V���0�����=��c;�9%�Q\�,t�^��S+��w��F���>�{��j���9v1��S�΢xU������fl��3CiA]��@�\��-+h����8]Ҧ;����zn�⯛�1$�]h�OTx�F%�������I�qZ�9d4�C�'����EJ=��R������Ȋ�����4���~�g�7�`�U��4�<���۱�����P�C>�/���]�O���������Gb<���	;��Է�-W*҄��V�s��������pD�(o�<2Eͩ�7�ը9���rPWZ�#tU3�D%umm���'Y�;^#����"S/���i�|gHFl&kBJ#�iX�w����%���ʲ1a���
�~=��7��<�׫��G�g\J��V�z�LD����i�<�5��~�q/�֗>�۠9}3�*:T[���;�|��bdS���=�N죭>Q����Y�C�1o?�0X����ye�����"Hq2�36e�+Z��_!K 
�m���*�KMsѳ�L�H$'y_7�QsK�T�Һ���/A�7�0X���?��2E�W�\�+��[��ω_���|ȗ�4����'ǥ�LU
���-l��w�?��x�=`��d�b�Iї��6#����`&�6w��T��ա���J4S�u�J��>4������c&��o���5Z�qg����U'���j�6J�����/%4�T����huġ��5�iT��p��O����T[Xó��n �udA{Iq����'h�������-� ,́	]��$РA���>*��%}��H�.^��o4]��Ov����v[l�-V��!�N(`�n&����;�ค���{�V6�Hg�S��$�A!�>��<@��Kw�\nʓ���2<#�=�0�V�\����+�s]M��������Y��=Yk]����8$ց[�� #� ;�|㪉�~���D���i=֭���J�p�m�}tv 8?�Q%^	�$&�SA�,�	)*�t@^뗫�iV�~����|Kq#GN����^-F�Q��B����]h���-`C�٢E���d(�P��]�[��������m`���GN�f\f/�3GR��%��|fn�Fa���y%�!��f����5��q{q��,�Z&�"�߲z^�(s��&���7��F*y�����U��g���@p	SБ˗�5U̴��OC�Z��^�3���8@�5��T`_y;4{�;�� ID���lMӖ>=��N�$�(Q�4���S��ı��b公2><��¶R�% ��(�mN8�E;�����,�<����������\��T��}[Q=xcV"ln��q���h4��+1�Ë��J�R�Sb�-�i��)a�<��`����������]p�"�=��y �?N|;m��^H��G�D�H���L���ƿ������r�Ek��/��o�v��>�O!�A��!h�.��^����Nu�I.��2jsq���c�:��u�g�/���Խo���?�b�:�H��s�A��`��E��rk�����D/���s%�v��
e�,��*�
�lWi��VLs�a�5|@�Q��A�.)�� Υ_�h^Q�1�B�0��N���:o���l�:*��
_�����W��H��r�fe���0��v�7��u^R�p�.���ɑK�V~{$1����8���:}Q�[nP����ͭ25��6�� ,�)E:�P�BM�V�.��>�1lC|�,��2�|����|�fs�����
���*� hHfX��u��vi���;/�6\�ZGT��ּ�K=RI�W��h� �`:��V	��ذ~a#��Ö6O��`=ؕ�藖;DO?	���`C�T��Eq(M���L`((�}v�r�C���yఊ�a<�8�eD[�CH%�@��1b}K�py=����lMV	LXE-����5�$9�F��#�P�Щ{��2~s�G-���E�r�n�i3Ss��k�{W�����MEтgM���������e�U�Ї���F������hk�Zi�G� M�K�����f@"��g:g�c��F7����Ɏ$w�ސ:5��"`L�B��'�=ԥC�WB��2���H n�+���y���s��G���J��� &����5�̽Dq>O�<��/Ų(��^
��d�pþ^xa(��,�|@<���C>���#�� WLe3�7b�T��>�r<o&�����uv0�m'�t{�}#����C��<{�'f�{���Yq������ێL�-oYx�l��e�������W�s4�S��ų�≹����kw��-�1��Do�"�H��	i/�K��˹�&�2`��Y;n��	�]i��]_W�����(Kv�Q�Ȥ�G9�{�څGI�	sz���)���À~*(.��]�ب;S/B�{ ���o���Jn��_]ay�Ly��Ci�%L���^G,�eFu���a��U�l��u{
lz�wt��sf;��}�~iX^�]܂įW޴S�����j2� �O�F���w`B�UVi�@���u�4 ��O�4l�U8M��\�^3}�r�J�D!�]���C��z�['��-�� J���R,�� ��jË���7�� ���g�
yd|5Y��e�/���q"��������������)���a���;�7��,�)xIE�����CҦ�wevZxgk]����H�ZU���Pgqr�m@a��,J�����H=4��D���G�g��j���%����w6�p� 7�`iv@�O�h>l�k�{�R�m=Ӡ�2my,ōR���"�(�B"~��B�T3_\7!Ra�kT�t�:��� �Gl�?nV��wx�f����V�o����9-AX��@������z���t԰pj�2�{|�;������ڣH������V.	<͐#��V٣(���yB��ӰP`�|6m�����1�6-��&!�K��Lflc���@���v���!\�QL����By&X'~��$gT�J�zZˡ������4M���$���8�t�8�+f���{,H�t�&�pU�=d�4�pH/�����K.=J��u��NPf7��q8`��qm}]ӹ��k�kC����� �����ے��M�?	n�p>��W���}��K+S�US�A!����8UZ��_}r����89�@Q�i�=���"39ބ���D3�p�� ��.�b�����B������YT�UO�K]cj�hӨEp?X׈j�1������a����c9�"�n��%�N��ۏ+'˗pp��;��{�I-9n��m7�SDʓ�!�`��1\ʺ��i}mD�όE<���w�x!-3&UR��HZ?�l5����(Y�\f�������@2Ħ�c�´��	����+
�]��N���.���&0��Gbv��u?t��8Y�Ϊ�^��*�]�ؽ����p�@�}:i"vo��N_Ϻ+Y �f��&�7n( Pb?���aL��
�/�S�xP�q�9��Z%�O/_��<��kRrUo��R���~�����7�d,�cn1I��c��d��a����f� #�zïz���Y�iL�1��X��0]�6['��3���/�����"���O�� Uk%B��ܛq��1��+��ɼ-S�����#��E9��,k��ĵ�^��"������[��� ����r�	��㙣z��x�}<ɈF\����j�%�V�
��C;q ��{�j{U�x�oFP�8�X<�R����|?�+�>�Xe��� ��h'�=,C���sKcwPHv#�P(��󀒋Z���U=e~������|�\����Vi��b���M`���:���+(bM,3�!�����`�3����&���~���Ǡ���&KT�8��r� s�РM���Ll&��s��!7cVRv��Y�س���X�q��w@II���h��\eD��SkU��_䧭ct�Q��������Xeh{�>n�Z�<5���o�㽜c��jR8?�����Qn��������
�3/&͟D��&�)��l�:��i֙�7�5|�����7����I���r�V0���)]/�2T?W�D�$/���7�*_�=�®��|����@�N��ή�m>+�������e�A���h/f9ea�l�(�Ʃ?�m5�15ʵ}�j�\k��Q�R���U�d�g�8m��@�T~����:�����%�&��ѭM���=
B��A�!��������A��i��NZ'B�/�؛O(v�Pz4M�<�C�[2f�C�=R�����V�PJ���`�L#gsn&Hנvț;Zၣ���Fr�{�����W�2�N-T�i��	�b��lK\6��x|��^Ǿn><�`Qb8JQ���XG�	�X\��^^n��3U��Q�,|@�W���R�?�L	���`������ۊm�d?6��w��e��R�i����U������\���1�����#NQ�������Pc]-o�9�o߆K��e�%m-�Y�p�V}����Zϥ�~�ǟ��V��	tA�m9eV<��'�w�͡ >�N���;㢅Q|�����;1A����� 3m L
��g�Z����y#)C@f�+{K��r�i���0�������[�.�7Ι-͂��?&e�7��d��h䙆��s??z`�Nfh�'2�1����R�3桤4��B�J�Q���f�dM��E�+n�^��&$������Q(M�[���O�@�~� �ɉ�dK��B�����`k���p�s�� 68g�f^�n�n[����T�w�XP�����@���R��M|`u�)-��l�,�\�(�p�Ma8A��@�����T�h�J�"C]�*��R�!�li�h֪9̨97Լ2���|V�c΅�����ÔJ��Hυ��7'���.22%&�YFl2#|*��H[@>8�j�J�4ƓvXlxV64EB    7aae    1400^�t��)cpAd�Q*�--�+;|E��7%.-���pDYO����1n�9��8�"��b0���d(�F������/(���AȘ�)X�c�<P�u���Z�rxl��
J�\Pd��Ӟ��T��bХ�
�^��q���F�B���*����ph02Ts�{�4tC��)���ɐc�Nw��Xn�>G& oє/w�ɉ�ϋ��	����_���V��'����^8tm��W�~8j
��r�*������-pj&l�Ԅ�.M�+>&�R�i�����ȴ����Ӛ����g��M��^H`}VYvTp��X�)�ֱ��_XC�)�ꝁ`���[V=���P�$���Zo����O��^�ձc�"3��K�\�S =o�?O��d֝�"����VWew�K�|A� 	��3�ت��/�ҵ���s��c��z�7y�� ӦS07עr�x�@$�y��#͠?��12���6�-z��v��v5����Y�E�26��oOo�U±PXD����Y���������y���\�I�g��\2\�k�xb�$��f�LK7�m���1v�� S�9m��w�����*�w^G��5\Dg坛��b��/ܤ|a@�#4о�T��h��5DC�'�=�o�����f<��N\qF��b���\[o���áh�=2m�j��V1W;��$�`��D�h��������[_�֓���жf�'ߏ)�ԛ�sl�w���24F� żs�JgAp�����N�3[���3!88�6Q�p�������z��ՙ�@���q�N�����������)5- H�&�#F��Σ2������7TJ��bY�RIn��MT�nQ6OTˣT�,*"$DuY���$�.0*P��W�~g���"	6�dU9��&�9Aյc䷃SC��V�� 罔VT���'J֓A�j�W!�"�s�0#�Z�f,��[̤�e�G�`�/7sޘ{LB/�.��5щ��[b�E��{�G�$�]�X�u���~_$�m���G��Y%��?m���X�����b,$�����3��O�I�9~�&��p��2�r�l�I8�sf�2˫��g	�?�R��U��L���P7N�1c��6�YXi������"y�f�d%�rZ{X�[���&���9=��m[�~Sx�m����4{�K��n�2�}2�}���"�O:�����5
�{,���D�.S��h�Q+:pC���r��<�Ё�#M�&ݢMp��{?�4����xC��e,=�v�e=�J�1��,PL�q�}o��iw)w
��w�	4\�,����l\8���p�e�8T:�Y�q��]H�[1i��Dk'���@�j#4��`~��-@d���d�����>Ɔ3ԓlG�8SE 9�Y���w=�|����:$��?����G�5��NޙRo��Ӡ��;pZ2av�g�'#)ȋ�A���ӊ"��/�Q��	���*�.�\W����_��T�?��=�$*zC���1kQnU�?<��+6 ������G�,L�%�tն�)s�a�1�f�������a��/Bʳ=�P8DJ�Ķ����܉��L ��H��M�t�Y�3�V̖v1d^Z-s�fQr���q����ؾ��zo��t�+*�u�bT��.-�tU�^���1c�!��p5�(-)�" s����uT5U�&\F�s�7��_�J�L��z��a׋��L$�>(�-*!7.�e�	�����/��tiQ�ܮ&*��vb�%-u���˄�@�/I��l+�"��?���wr�L�t�U5�lo(��{�q@�����A�0�YN^*N��,�����V�9�qs�0D۫��F��E�܃&����>]���+��lPR��������?`��|_�6`w�S���VD�E �D:�ąl��j���|����{JڮTc��D�_/h��7��1��P<��~���g�>;�����J��$��M�U_k�����)-������L�r;�L�;�`N��NPLÊ��U�{r��Y�ӏO���]22�z�P����h�� qd�G��{	l���&���uc�k(sXN�=�� ��o~�. 5쌞�	��S~���uX���]/CⰃ���S�v3%��)���/ N�����؀�c�B.���9��[�`�0�5��p��R�E�@.`������o>�w	u���cCl����	":e	|r�,UhC&���PD#�siȨ�?�jNj`m�^r�}�����0�A����C&���,X�N�_&H��51҉oM�zc�p����{	�P56_�?��~+qKÀ	LX� ʎ��#F���U�O�9ў��sjE��oD�st��I 7dDe��gP�rǍ�w,���yb��+��<Q;[��M^)� I!'f��>czf���fO�6�/mˈ���s%�̶F�O��:�=H�3d.*rd���u�oh-##Q�b�F��0�d���
�����1D^�\�7��w ��Y���Er����c�CNDדܾ��ͮ8ȫI��D�����~�M��"4)5}����Yg}|��6*�n��-ڱF�0���*����yX���,mnc�'g���'T����-��g�V�ZA@B5��.p�CJ)���o,CE��������ŎF���k�'sO��J��ا�����R��*w�_�.,t���I�u��u�o����
���H��t�vB�v7��4�����I܃�*����C!y�p�Lt�����i��H	[�΃��%��A���~f@W *n��؅�"��rBm���CP�FL�-tlC�듿=�`�1���ʬa��{vX&�4��}U+�m���5�Rg�Aj����X��d��z��2�0�un���9�i��B�N�p��F�qL3�8H�uv/
��7�v�rBU���1�P��P�\��+�gK
�iP� �(ո���<���M#"1!*����SV��)�{�����A�j���\��]��|j��O���m����o�s�Ôֱ�DS�t\"����?�(Mړ�>�����+�.ǰ�oR|2`䮗Wg��˫��ⳣ�������:���9:�r#�/�]9rє���s��$'�����K��!�;���p]�-^��(��c
���@N�q#�l�6W"�/�q���ò.e����&�!x+�ٟ(j�i͖�%z�[��7��$F=�������L+�gX͏�0�8h65!˦� ���M�� ��|��<��B�3R5�r�s2�crE*%N��x|�v�;��x;���JGk@�=ҷ��k����Y��Q�*^��$qJ�� h��L𙤂�հ)sE&�d`��a�ԳsUÖ8ڲxG*U)����R���vR�x�9��?&����w�����s�+�S�a
ܣn�L��A�K{��څ��n�k!T�c�����H��_�
5JoP��ʑ���7�B���t���E�FO����h���x����Uփ�)!2�N��	��_�:��J�[oF}�St�@�t�J$����#J�#��lW��JI�E�ʞ�6��/�'ML�XwOX��"0����Z��J�1�4 +y[����x)�֑�n�,��6���L�l�O�Ί^ZDk�w���5Я�<0�C�$�ٵj���7�Xta�1��^�󾒏G��jz w�of#�p�Z��eu}s��_���uZ��}K��5��O��QT�y�vo�C9dQg:%Q5#Ŗ�ֵ�揁hܑ3OE�)a��.�m���z�OYO�=�3Y�VhѺ�I��_�u�j�*+�}�O�ȭ�b���!��7G^�����G�r�L���`�<E��9�$�e�2$�[�.@z����A�mOoD*��X��K~�� |���T:#���,��lu1��X�w�=���F�� ���S��	֨��X)�d�u�p��&أ��`��8�Ҫ��Q���s=y���`�Z����x3�hEm�dC{�<}�_�u,n���l*Q�")��#Yn.z{h�j>�<�c8sok�� �Q&� ��߽�<�q��������x�6N�}jկ+�
|t�x&�;��>��~㞮�j�B!�2�*}�z��T���N��ױgIt
~�����#��N��yo��8|bZ�Ǥ2\rF��Cy�;HX�\�%N�ɇR8��;��oƬq�qN�t�G�WG2�ߪ�2>�!��(���XC>8K�'��Y�e�|���ڨ��v+�Ϙ�A7ruLo1��X�a"�m6��}�#���A���0��n�rI�E/��3���8}�3�Ɏ猍�#��ަv(m���"D[9�}���#������X�z�Z�
"5e��<�i�^���ji�xi��ɪ㠪u��A�8XT7T�4��&v�PS"bf�0�߃8\皹ߤ����^SB����������+A:���nN�m&��>�"�x�\�4�ϱ�V��Z󮚑�6/�z,�L�g��йI�?��<�����L�����"��&�:K�1��n����n�<{��䙘���ˋN�V��R[At1�|g�o�i�>:������!_�!0��pݝi"�C���8(��T)�����Vy0욃Y���(7�ץp�*�����[#�U����:#ϗ�.��EK���d�%����Ų֩�~�xF�������w�wj�����}�V�c�@�X���"��}jY��B+�z0�st�m�B�=Xh�Maf�:��HR��S��7�P$/zZ�a�BLnX�.�_��`�U'�U����t�kKjn���.�"_����A���ϕ[�q�	�9��z\1a�Gﰄ$�$�;m}�դ7�( 3��Xæ����>��s���zU�*b�qɊ���ȳMӱ}}'0-���w�TB��[�φ��������uf�q&b��'����6L�gsd�!����LkI�"�2�<�������@F��t�[���޳o7��/�������z�����"����6�x�C�:S�v�
���㪡v�y`Aʉw�쨁��t����9̇E]���9LN0�;��