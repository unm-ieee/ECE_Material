XlxV64EB    fa00    1ba0mHb�%�H�[�A:X�xn ��@Pp�����k��4g��F�[\o��=��i:�3��7N��ԭ���+痠�6�vq��S��WT�����`uRf�[$=��C�J��ٍ����;9�-���s#�m���}{X�xh�h�B0��&�I�>=M��/���=���l����Ʈ:�:2rGO�!�H�_��!PtN���{kJ�b�F]T�"r� ���fL)��J�0l���>�O�b�D�r�yB�en�)����?M~NACY0qG�N�`�"W�Ut�k�(,��{������k�+�W^?�W7�]���G�ӷ��=6r�/��s��`���.�`����18v�OA�2��Zr��f0�T��.u�2��<�:��κ��w�<b����g_�m�::���v�Ԅ��m9�z��"���J�-D`�EʤIC�s�H�����ы�?>��~搸���Gq/������G�S���r�'ԥI�ǽґ�v��#��]?݊�~izeg�g�Y�]�Ma}*od�-Qs4���$��$�2�t5(]�n'F�w�y��s��q�ɄB�-��3a78���V}G�[o�W�	�=4m�?���y�29�u�ܜ<�����^=�m�:˰~)�*O~w\�<~?t��A;�&�����J:�r���d����6�>q!C��pQ���>����+����ŅD�c�L���kE���X%+��7r&��:5#�_8."j�����Y~ǮÃ# ��9¶�����u��j�C��75[�vj�D��h����A|�7�)S�T�
��"agݧ4ne�<P�o�?��O�^���~+��í�NN�����F��\�v~$Ld@ʬ`�+�6	�&�����
�����Q��W�Eb%�P��h�.�Pv���?Q`¯,������6�]���+�"	�M.av�������\29A�6asi����4���$�	BP��v|6a0�	�G�� �w�qG^a��i'���f�&���#r#�^�EK�Ka��,0}�b[���2(Hl�6.��&v,�ƃ������S9߃�GdN�q���)J����p 9�I<�)U�]�Z>e;�)�{��md'��}���~�g��r���f ��)�������늰!4�WJn�
��U��L��e����';Q��3�e;T~3���1�I�����o�p�8�raǬ���7�U L#��*��+��O;�
�n��-V� C�,���3|�ՙ��&�?�h�y7=��<�zf���@��X��0��C�J��j�8ʼ�Qhg�n��,�P��~+����q�0%�a�W��e7�w��kj����.��r�����ӧ���3���fusI�����wm�O3]�����;��E� ��R��U�/.��6�`+-u�0u�^(�����|o���S�U	�����@݉_��fE��Q��q�
k��r�RX����d
]��ѐp|���2<�|'�_�k7C���� �	��;��q�����0z|�������oW��6�.�{Bc]�����1#��,[n޷6��4}ef�g{PSbo+g\a�a%%�jQ<�}�/�f�� 	@�m7�VZr\k��� �wS:��.,��q�>�WCh�{咏�� �����乺j߆�t+���y�U'�g�f�I솳�`�+l"K
��k�Sz�)]�x�d-�$(!���ذ��T��<��QñNhâ��B��
�+k��&�"�쑮:��R�w"duJ&���b�Z�ً�HE��J߸,0�y�.���xd~p*j~�0�=���.��e��y�M��1W���S5��������;�yd�hB��(fA��j���	��J���[h��gQ
������3�Vw9s�ׄ&�<7l�����[p��f�]�8�]�;�w��0񎔴A�*o�24p�V� sx����Fi��.e�9�G��9�l�@K�<��Gt
A�	���EY���ἡG�_K~��cJ`���ɶi������r���(�L�2d�]�S��������y�lsҰY�#�a�^��'u��s����о���Kf/E[Ԁ��"1��:8��c�5
U��	�^Q����9�K�e?�Sl|��}�˼�7�ż
�P�^�h��Nf*�"c��\ �a�����D*�Y=��i����J6�3�A��o��k6Z�<�y�ҶL�s7�hS�Xw��AnzQH;u����vf<P�w��7�tz����Sߪ�3�˃��qL�>=�`Q�,a��a*E��O�]GG�3y��kA�.�@	%3��["W��w~�2���bN�S~�GΑ��h�����0u��Lla]�S ���,X�`t	@��i*Eq�t��y�ǔ������&�p��U *4}��ɋ0�b9&�J��:�g�*S��9�9�Q�ފ��C)	�C/�K5EF�?��b�9f�X�|���#�g����P����pˇ��qߌ��"ԅ��dR����D���T���dj�9v?����נ���c#$ց)�(	��]	:{+��u��g0$&L���K
��1Tw#��%��6�Tw	�ʰO��H�=-���~d�_,����Z����i�(z� 2Q0g"�������;hR@_,)�8>f/F�����YF�A1���:
��}��u��C�������j L��q��c�/�I2��=n??,w�L"8Q
2���`Ɖ!��r���_˨V��'`�9��e�)�?^�G)i�+��|����M\9�Γ�C��5�.4����΋��ݕ���c����P y9�gS`��v���-���W`����9D���^���vN/x����+��g�v�5b�ޱ�:[yy�n���4���N�z��"�x�����}�N�H��T~~�I]��F��f�@Ic|zV��3���{����qrG*�O+4z��ՉɨN��EZ1�`8/��t}�1g��ɧ�󯃿�?|:n���;�H���yZ4�ה��7�Į�T�ƶ�\����'�^����gp��U'��a��J�f�Ĉ�\�!���4+sKm�q��
���Ri5VWō!o=U=���Š���ߥ2ƌQrHxR���=g#���v�3=�ƍR���Q A�O��W�#�<t����?C/ɂO��(BF�Z��;�l(��B�98�[���@[7��[����� /{�!�	QU�"鵹|I ʭ����TҔj��''�a���̰r/����{��7rA��!��m�F���y�T���
EI?��#�e�}=<�k��ͶOr� �8��8pW�6��S	��VC�]��6��O8��;Qt��Z����GO.�A����̬S^[��f$s@qǑZ@M�riԎ18���Ԉ�8�v�X�����B�Un��ݘb�Yr������M��X���k�<.�+Kn�p�0�hd��ᤰfE�T
å�C�g>O��,"
�ӠU=p����VUpБڿL"޵��R�fW�X�=h���u��_.���&�����T�8V���6�Ң��/�z_���ƅ����e��r���dprEiFl��H�0�l@P��_�riǔ��(�BO8�s���Q��3M�{L@����l$NS�5��D�C�őR��9�)��ܡ�8�j^^Q�:�-��\��A�r��ty&���lAe!v�,Om(=x�'�D�	��">:k��:���a�w�^N�a�n�IY�o�"��Q�30R{
-�드o���7��Jj:R�U���F��Q�������4g��q��V�d~�4 �q���$�Xo��P��E=(v�*J��q��'��(o�٣*��G��wq�����uʨ�|H͠��N�7���s*Dyo*�)ɷ����)��j���_ʔ�j���_E��UK��P�:�KU�O��iYG�`�g���j�T7Qz���e��l���>��<�0��ڟ<��{�VR븾���3g��~�<=X���Qb&��g2V7����Ĳ>@���r̾T�� a�4���?o]č�������^����&*'����ƈ���y�م5���y��Z��I)�qX8�1�)K���l��?�7u��7v�Ӿ��'^�0�@�[<A?|������$6B(��� ��?�b#�C�R�D�E>݊e�a�y�C�H� ���7���AW���	��5Dw<� ���vWQR?� o�/��>6F?���x�qt��FmowT�j�o$��'��$�]M-��c�HX��Rz의#��#f�|�g���ָ�u'p������]���@�� g���;AN�
D��
���ZW�j&n�R�)<M�O���\���ӰqT�gA����c x�n�C�nNDE���0h������Wl��]�<,.昊#U��dY 9&������ �G+�/�S�*v5���"O$Ď�~e�#lʙ��_�|g����	����U�
e��a�GR�I� �5Q���g��3�= ���V
� Vў�\���Sid����NP��n7SBX��u�'�UW���8�V���X�+G����-o�Phyj��+��_�p�^�2w�A���	0ϲ���:��.'���;���w�"6���T:�5���-����i�4}����x��Pw�@0e��dW�]��aiג�������7u�u)p�.��.��m�e�\�<�9�5xA��h��y�K��݈FT,����h��z|$H��.xCe���\�N�A_�ќ���&-��h�(A?����
(��]*�6g��k�U�h�_����U�5>8c@V���/��7����Ck�}�z����;���?�u�w"j���2
#�.�=��ڲ�p���XV�V�>���OEy�y����K|�$JF�\N���1G�hv���O6z��ۂ��J�o}�:�d����Z�v�Oh�~���n?Wó�Sw���ŇCO�~,{�u���d�lV��H���AF�u�E�W�N�L4�T��p:�Hs�$��A����?PݺH,�q���u��:�=9t����`h����Fg�X�*���AY*x��x�@�ݜ�a���S�j�Tj��n��S�l�!e"z�|��u-���0�{'���8׉HWDG`U;hW*D!��Ʀ�t���/���/��=h�7�H&d�Ik�j��=A�ܫ�"-h+�j�R[N��i��wEԯ.��)_��'�a���*u
&��ڗlwo�*�G|[�O)�[� e���bg���]��Wq./�<��u��FJ=���NP�a���6��(��XmĕduDhc!��ˌ�<G	�K�c;@�irF*�"�4�1��d���Sld�����4�b{�[����ݙ �+rw�~�~뻿�I��wP�inE&]��/��W#�C?��5k4Q#
ײ|���Uswz%���[�Ш���21�V�0)ª��pm�>v��#Tl����JW2"{��'�z�D��vR�h�p/�V���ǚ;伜�/�r,� �ջ��aNb��+�|dE�p�����<�����D+u�_�uP������c�&)W��uFt�"�{~$�{hs^b,�*h�x�)�~��"k��x������� �g+�Q�	���F��|���Ld��\���s±���0��L?	A�)ｫ2�m�*DW[��v�t��v��Ρ�J�+��\���d��Ʊ�ό��>�ujnJv'�{`]g?��"k>�Z�C�CQ�D�7H/��_`��c�)�9�fd���-��$Ew�{&Ώ�\��ګu��KW��<2��m0w'Y!"�;�%���׺�8T�!�:�^�}c���.�j�A���f#�{�?ˇ�k��B�	�:�������wn�d(��K�C�����@ױ}��$����nx���՜	+��-!�id��˟ҽ���_���G�W=��{PS���;��I���O/C��jr׷^G�q@ۈqq:o�ݘu��=��m�m�:���w�@������2��K��k5�I\.�����:�PJpF"��m�n����^"�? n����
P�����U�f|��
���L!��;^{�^��)�7�>Đ�dnn��\ge�Y��1��6����;�{��dr�^��U�DB�pGk]u �"u"s(�~j����ɑ�̱/'c*��n{pz��4��Ùy\�^����fǿ"��y��v~lFFBWR
	8�S�x	:���x���5($W����� ��Y��y͛���N�,�G+r��3<�g�L�?��ô�D��x��{B~�
�����q6Dmװ�J�0�aRO�	�#Ź�ha�3~���C�z��n��I,>ZpvIz�<��F�xz"y�ח#�U�:@d��?�>���D���s�I�2y2�ކ)�L�z/��^+��nk�T^�8��y�s�v�uH5 �Q�64f� ���!�����e��R��1�+�y������6��v�S�r��&�2eCE�6�5?E�y�����1�w�:�Q�0%����FXl	7#Y?���*?�{�o
T���"솨�Y�@c.�XO�l*K�VM�G�sCe�66�W�v�Vxd��������}ȥ����pdڜ'��W�'���=\=$h��΁���P0�$�"(���K#^�	h�Q7}#�va)�m���L�1��A�z%=�o�uk����n&�P���B����@ˡ6Vfә��wɮ@b�>8B�]EY$�� U��(S��zz&U���"��oj��Mrh7�b� �W�!�ʕ@3�6*��ҥX�%�s�����!�Y�8 �j�'�*[�lcі�s�X��h9e�ߚ,;v}\bI�<nAN�"}�,(�Ց���i���n6(�*�%���?w�g!� n��:@?��]�LB�=@�Gf7��I�'��"���i �k�p�py�{�y�˚e�_���?�Ů�c����H��²�O��K��
�����G���Ҵik�XlxV64EB    fa00    11f0!��n��A� ���$z��wV�g6Ӟl���#��L8��qv�h���}��!���j��CZ�i��	�O���W�=�Y6���[�/^*
�-1�� ҫ_}�������@fd���Ky�Y`��L�z����p,��+�7~3�BI͙B[��J��Aw��U�^�H�4�߉����3����{m�=U��5�O>�^z�F��xv_`ǢQd0���>�M|��yH/xyp�n��Tm2	"%��n�#����h驮����3#�Y�n�:�h�jD2DC����d���� sJu�'J����*e5O�	�b��I����C��H~�01| Ad�4ba�x_�6����`�W}�v���Rs�d���fA�"|8���`G�5=�&5�`��ᵜ�ڙ��O/��x����wJ�VR��7�kV��N����Z�f���s��?T-�2��$����{�x��ApҼ�J���D)�c�G��R���T�	7j���h�6򶕒�%�������&a��������^��y|�5Mֳ���^�^D�/f��W�Rb����0�E�}#TMJYvz�g�3�_�<�uf�Y��d?H�V��+��gਖ�f�3�W�>�K3���Q�m���3QC��0���0b3�'�#xC�AY
�z�B�a �x�(J���ޓO�k�h���|F��x��;��ydVg^����\���/Ɏ��=G�R3+�����i�@�����J/G���ޤ[X�0�N���m��a�z��h>ѧ�Q��xW�؀~V�	ovd�ҏǗ7��6Z\y},c%e,�/��K����I&4޴'�\�9H��� ]���Y�,�2kU��|��|�I�B��ɲn�uŰ?9��r��]wY��^�U���	w��U����ƍ>O����X�������e�	^7}�-�F���4u4�ᒶ�n��
"��s�6�n�#�TU���j��K��Cm�<i*��6Г�1� LD�Ny�Ɋ'?����;O���[Cf��+����$��H��v���$R�/��fMl/N�N/�n�	���z�4���=5
�yC��fZ�R����-�Pn�]��	���s�Ug�u��>z��f���ѝ��C5pHe[�]��
�z�2��U���'���Q钯v ��Ȩ-ͰG�b��ĺ�lM��w��n�䉻jX���� �>��9��X��v���RK-��2U,�_�)�#�if�<�>�<��*����Z,�"̚�0���McC�hQ��q͊�#�+��MJύ��DR�|e��R�ւ����C�FRzSoL�@��!^�z�$ѣ�0�!M�j�5�� ��B���4N�"�@�ޏ��A��+�Ζ��*�Gٲ�.���F;r����&��o��V�~���ϤM��4�;ײ�B,������{O�]�B>r���g֬q��x�Eb��+S�R��Z����/��&�M����#2���u��A���^�����0�g~���&�ř�\�6��4nA@�Ұ����䘭�|?�,�tD���#���@�9�v���z��ٟ*jܝ<h�}ˀ���>'��_�qq��p$�U���UB�����9`jB���擛K��3#�v��@�J|��ל����k�s�f�5�uz�F>М�(@'���!�i�Q���˝YͰ^�N5Ѵ���~�#FE�Mh�k�3����bH�Eb&}Ĵ37�g��r�{���jI��t�0>Qx-/�&�O/]�_���,�grߠ�٤��Ӝ}��x�XHH�I
s�K��Ex�~��R �U@�tК��Į�l����K��ͬ�K��O�	��V�������Ǖ�m�$4`L�7C�9��g��f��f���׸�_�qhWn��#�c	^�5]gS��nh���kv���+C����7�n�lގ��$+zU.?9aƠ;����5�Ӫq��ޡ�v雗cEi�Tmhc���I��g||�ͭ�����گ��ʙa���X����P�Վ��>�l�(�8��y� \�@�:��9���X��<�*2
�k�~6!,F����H7~Q���+X����Q^���o��N2�������^�q��q]I�t�V�N�-�_b���i�IAg��#?��y�!�}I-��|p��8Py��x��I�� >�4.[�Z�"N>+��i�l�wبP^�A�I��_h��n�����dld@M�.������x��
���e��a�^�,�Y���B����z��=���mU7>g�U�]˥��ȹ!6��B�5�ᣓɼ�� Er�a�=�T.ޢQ^��ǫ�ٜ�fb�J�uS8-����>E�j�Wդ�q�Bi�����m�e�Y2�����ܦNz�#�w�N xc b�m,�ȟ�	�R<#
�xu��j��dezf��;os��ԥ����H�6�0�F����۽]��2��I�1r�)m�:�^|��*�7���Y��@�-������A�EdW` �MAȟ䏯�:0g^���y�A��Ѱ?L*<�zVY��Ʌ��*���Պj�J+��n��B��I9����F�`B�I)���z�:'�:�$G���װ~F���5��6�h �zj�B�\���������XN��+�Ѡ��R	x��G'�l=و���O�b��R�,�[�3��O=�ԯh�D\@��.�{3-�>3i	Ë�N���z��c��A��n�3I�qxx�6ә+�\�Kn��zC�i�a��d�L�����*��$���9!dRUe��!��9��zUOWi��X��s	p�ɛ��)3��R�l���]<_o��T�us��et���	}dd����&@��#�N�GX�b��]=W�D����*���Y@o����l��P�:_�_�(WϏ�\�w�����jp����̪-aK��J귗9�m/�1O���I��C���f���T���o�.3NLY�QX�.H�/��%7��X��e܀�S�A��N�>���U��м��GC[�RLhеxal�[q��6ʻU�w�Im$�9�Z�V>�
�iZ�r���3!8���m]G/��J��rWo�<fIo�o��s��k���8_�j�%o����E0�������>��c�N�|�Zi";ş7t�([�ń�۹��!�|BY}i���b����`p�Ѯ��H��x ��h��0d�tה� ��
HҊ�J�c��t'�-�:��݊���iMYt��6 �<�\[Ǒ�XqSåχQ��!]Z��q�ui�K�i�����z�"ć{��gƯB�엏{\����	D�Mۑa�R� �K��]G��G|�vqUm���#�"T�e�*��2�(44�ݾ#��/#��p��j	��A�W%M�ԝ`�6}�.ܽ�r�/ �J���,,�'y�"� ���]/ ��/��6��b��*�}�]�Ш���3����U���q�Y��R��^J�<�N��J�9+[D�m��햍�q����Hk�m6ō�Ӏ�:�

y����b�2���Sg�pdF�)������h��m@����ނ!sg;!�d�T�h������F����2�SNj;O\Z��5D�fv����
��k��]u4�Tf�8R��z�tH�Tn�r_�
X"ec�U��D�;��������$f����B��jQ�N�*ێ�TSu���c���nP�����N�0T����
�1����Zm���&)r5��5c��j��b��U�6GcZm�HF4�T��� ��t:���[*C~X����ݠt.]~���ܿ
( Ϸ4�t����[��Vd���7�ȟ��������J�7#`�yH����ך�~;��yI���t��~s�;y!��/(�e^�D�R�F^�JA@��Q|������'6+Xg��h�8r�����I�g�0�v��+��Vh�����@�%X�l���o�$ی�v �[�z�2�J��L��GɆ��/'�j�3*Ϫ��$]�5<:r1��s���}��=�!AVD����;v����j����c͕֮�6m�IK�4���/ex,
��JD�à� h��`��sᵨw��@���֡��`�`<�P���������]�x5$-<��F���mo�;��#���gE��syYQ�r�q�
#�ֈ�UN[y��܊4�f���B�e�@{�h7�� ?����M��gJ$-5����q�FK����sj�~�&�'E>f�L�<�m"[�%=�������=ō�P0p�xa�M~�
����?�\z"h�H�m[�t� �;rd�A�-{�>	�GB6*=���l�i�\���SI{g� �R��T�ܡ��6ۙ�$�}?��|��?��!l�5��o������Ϗ�Qm��T#H���
��p#����I���"P�҄�߳�m��vF�(+[vUN�!����	��RB ��g1|V.��5��V��]W��"I`��Ti��	}�vU�lm�y��辬Z�i�
sǻm��l������Y��c@�G�r����E5Q7�ȼ��D��X��Ѭ��,XlxV64EB    fa00     7f0���K����g���9�e��B�vL+���S�G�����B�h�[w<������4���a�4p8<ֻ����J��d��{�:�5o���Gv,�b�~�d�P	9XP��c(^ C |#m%��Nw��/<�=��RR��k�;oc^Qq�Ӆ�	�3�ەq:�����욤:�%��;�Kx�%�����`�"��u�S6V˞� հ�Z��J���Y���b�'"osٸ�%���E�p�+�c.	[*��!�O9�A8�]��lX�����*�/�8�D��<���f$]hR�����sҋ
����{2�3I<��.���z���!��k	b�	S�ȌеV_���Q�u&�e�(��~ ��x�e� ���N#B���o1�`JU����KAֲ�uU�������O��,�����4�7��cW"�R�Q��p.���cF���J��ߠ����r^�).ε9��`fŎv�����"X�vIc��HS��.`�t�$����|h�77 �CƼ;7G�� ����-�����~�A�V�%�ǵ���[*�k��v)��;��;>RjD-�o>4vr�����gyS!��5�ň`���y �@ב��~��j�3�gr�ޯ��]?��l���Z���G��V+[�jJ��}%���{~�Q��{�ЫÎ���ۡ�jy�B|v�k��H{9�!j}�1�A��/�T&���׊�I�E/�p��G�j�¿mUZr:�翫��b~��m�Mċ��1j���.��_�P�T�C��`U���_� �>�����.]YFM��`�R)@�m����������`��&ř�I t"�Ȓ��"~t�1�k?-葼�+����֔-q��j�����X�{]��
~-�߯|T�@B� ؇�"=�P����s����� _9Ȋ,,��7[���<oi�����o�E &�U�]*Ƽ�x��8�m�P5�5��E��$v=�)��p&V�iy��9��>h� q�1�ë1��/揨@Ld9�(�A��.���;=�ޝ�l�y�rd�E�L�_�4�;�0*����Mn�Ru�@.��e�#C&�+���$���Iʑ#Jij�%�	�����xZ�*l��\��mw�	���r�ş���z�]�Յ����{�� �����[-�j���7�P�<�$΃W��ok�n��+y�L?O`�Z�i}/��X�$�	J�4��S��A�d�z��O�f;C�W��`I�hu�#������К%�B��klq��t���)��d�x�=�# ������H']�4F�p>�]b��>̊�BYhA^n#\�oq�B�I���m�n�����+O�c�67���e���vˌvB��
Kd�W�n*�����[�zq��,U	�ɛ�Ğ�(8�������Q`�n�k�qr��ek�m��4����BD��vvf� =dN9�W֤nf�79���6�2�(��W�����۶Z�/v-|��R�xe���mJOf�#_٩Q�����^|>֞_WCW��8RB�R5d�"WZT�-���X����Z��u��\���A&�����u�'�tt��k�#H��Yo�S��ލ�H��<�q�ۄ͑Sn�H���)�.�ٲs�㐚M'��X,7�T�m����@������p(<r���w@����?9��!pR��V�g�]�z�X��G 2�T�o�{�(O8�!�+�8$�S��䣳lw��� o�&tG="h��S ��	�z��s������B9�L-2�j�$��b��a��_���#�RFV�W�_1���A&�rk�|����9{����~L�#W>�����z����kUU���?��ӂÎ�;a%����1$Ydp3ca(��6=3Ks���x��O��
ZK�������ez�ӳ�!���A����nl����W�i�O����cߨ�p<�-vw���z��ډ�n�k�]Q���vo� �lB���P��V㋈Fv\�zK�ƶRI��|õ�XlxV64EB    fa00     870G�U��L�x�Yb��k�������P8p��X�O��5Ԉ/4#�qY��
�P�M�!w�b�e�Ur�9�J��w���u�'I���8:�X0�vL�CD�jm?�r��f߮n�By�5#H�b�W$p�-�q�����E`�au�q_sy�GH����*_��
 �l)��L�ul�+�?�!��E`�����.O�%�"0A���T{��A�w>xv��5)�"�`�)*ګ{
7PS�kV��C_�����ig;u���R���SS@���UF�nդy�|a��>��h��ťY�S��l�l�O��+������й�>�.٧��M�_Y���iy��Js���[��2o��.�#�&��蚌�.�п���)���?���6H_<E�dVrrP��{W�+�y,�\D�/�3y�3lW0U>x创YfQ_.�,E����~�16��r5�xmA��PBm�\.�O��s0R���8��1�$f�ȿ�œ�dQl0q�7��u]�0�A�γsH�rtz����:�E�����~�za����[T娜��;��r'���+ρ��-I2j?��u�L�+Y08%Q����x}��i:�붵%�l���Ä��N<�ع��>�j�a����p����� l��ሠOU��p�NY���L�dnd�[u�-�C�%0�e��$����I&r&��^S���U��p��\뀺̱p!ߣ�R Wp�M�-C�^D�J���D9��<��b;���(/�NX����ie�I* ��%N�>�r���	<�i�i�5�BqgRbh���R��?�m5��!=�I���8n�B~d �e� N�E�5����Īf� @&?�,e�'N��)
)=���F��}�_��{>��P�pVEZ�.�����p�-��@r����?����6�G���1�]��f�em��B~O�(T�~!�^�\��= �|?���;���H3�0�9^W��S�fo��t����D�ɪ�4W���U���Wr%a��K���[�@
�����-�#��`Z}�'��2Ҩ���4�lC�7����8NK��h�<�"�,�A�ػ5p��Ҥ��C�ܖ���"��sU�����:��Ӏ2	����|.1fS��H��;X�s��']��+�jC+�h����@D$��U�����p!�N�g?oN��PCß�1�.ݿ��J����`Q�r�cB*��N,�>2T6j���N!�9��e�c5h��9�1um��sz) �&z�wwm=�Ý�@�i``��2`�[X�I{��)hԲ#�̓D�?23`�,�ӿ5�O�D��64��V�DV�a�̓�Nf���dv=�|��.������/gi��a�{�q����Q�ݛ}�B2��h���0A�T�u�D�@�������1�pA��Ɓ�!��y�\����]�F�T�'�du�8��(7ͼm���y�Ǥִ�sG�ͥ�Z�W&%����[^8Q�O0Q�.���9Ls��v7�i�z����\o�5.�z�u�9+ H���!ȷ�{0���T�^V?�Q��w��x�lՓ ��P&�K���#�>%��V��;��]U��CЀ�&��b���{ (9]ʭx/�tD��'p=���.^�e�|�B"���ɫ,uM�TzР똊L�6���O1���@�W��Co5��F���ǟ�#NpqeB��k^B�����K��>�ׇ�#/�����-�K�c���k�u���8o�k�[�1�Ytִ��+<b�H=��"�,�U���[ѧ��{aZ�R$��F ���b����ny�!��lkh�&4������Ԕ���),VBJG%r�w9�4E$8�ϏWje� Ѡb'�,�p'V�N&�(ь�p�G�Ms8�Ղ_�!��063�R��,�ݐ%���5�Y@�4p��jAnL&�ő"Vm���@#���霾1kI�(��]m-�E<�Ya�F�uZM��ƣ:�vq1W97�Ű%����"��QN��t��J]�[;0��s,��Y*\�B��KjQ���)���D�8liC���E��u��л��)��l$:,9��i�[y9�Kө��Q	+`?<[ͦ	%�x9�-neBԸB�{ ���!֖�`�6�u���XlxV64EB    fa00     4c0���zE���_h��A����L?V��:&(P���3��
��瓃�k���p��w ��@���}�g�S�c�z��'h?n��C%�.�����F=�u�
@�Tc�3?�xB�d1�u����u���p�Wq��t�`�3�|��9KqA���m6�ڴD��0���saF�aU��r�!'����;-�ؾ`�7�α�G���Z���J$�	"�(E�ˆ�x�)��g��M����0�`�N�Hvܶ�<��d���$%�F_?4�.[�eL �M�D�y=L���f���[&�^���S���z)�+�ِx${���oμ[���QP7��-Q8kp�V��ʪk�ao��}_�o�*���UE��>�~%>�z�4L����ij��J!;k���S
�3�����`e��a�/�7��s�����Q��
[�C���g�?����c؄s��8r�zG���d�� ���^AXSF�Fbo�ut��p�))�O��d��6���
'6��A*U���ؒ��}��sod^PDk��Ԭr�Jk�3!
nzL������;)��Nto����v`0yo��xn�wi ߫������6��u�P��
���I]� ����6��_)��I)n�u�q �C�3I#]�`f���"v�Y0ӿ���|�2�+'F��e���Eػ\�+Db�8�7	�Xq�t���E�B�5�/8��u��=<�����tNr�;�P��׏����ɶD,^3AK5�HnG5'w?���]i���
������I�:��gL�$7����΁�w�	�yy\C��>�݀\+B"���@>%����债bG�2�5������CLňk:�C�n��Y?%nˏ����6r��Sqh��c�
ҧei8IC�acN�?9�gG歡c+JH�E�L��O;�=�)Nt���M�MfZ�OB�X��ly���ZF[ �<%�)e����{j �?�d�'��u���o����k>�����c!n�	H �hymBv0�!�M�҂�L�">P��������X�����4��&l�ӿ��/�v��i���OT����>��\�r��$O���bE��<��a���ɢ�T�{��s6�n��,'h9��qȶ<ţ�7��R��1�Q�L0�X���X�Vh��q��	~��g���&��
�q�0ڴ���O��">�+�}xX�I�A��V�c�Ζ����XlxV64EB    fa00     5a0NDv�%J.nѲ���X{�>%���|$H5�P���tU8Y	���ּ B�#9�3&���ggA{޶[��t�0����%a��?RnS�a��Ɓ��"�p�� jU5h��-�������|�M���?���s��!�$�J�(Meӱ�s	fq%iTL\������굥u�ߑ������ +�Q��0����l�l߮��d��a�'��"�f93|��TT&Le��-RU@�*!�WCwP��K;򉲙4IeS��g���)e�/_�N��޷ ��k~*�k�f��߂�%���gH��sn�"0"��&��D�P���n�ʖ��HԖć�Kto�{N�&��6�4�O+��˰Mڠ��6!t���*ҧ 3Қ�S��[ܒ&�pr��p����c���LG"����p�D)T���;�����ɡ�/[Ш�� ]5o�\1�W��N,�����cKg>P��t��B��Z��y�.������=��$�$j>ae6���lf������L�3���T�j���K(�s��IF���)��.e|�U~[�"�J.��:8�Jy�g�>���7��D�A}5��z+�^����2�PJ'9?��eg����1�J�����J���	�=�5n�|��2�0���E5k_�:�?�v{��FL�8eDD�!�6�X��^�P��(�<M�#��b٪��\��N��Z��W�M�FÔB�y��2������U$�j�:W�u��0���HY0� ���:����5�~��%O@}����M[��m=��-��
��Ig:�oT�΁3I
�m�mA��� y�۟{3���BQ�`z(���,%O�ù[^S:Sgj��Z��(��������G�m�!����+���G:Y�{ë��t�x~dzw-$`	�}�7�$��`e8
����0�+������¸>��@--�p��7��T�)!*���BB��ƮZ��rݱ�2wt˶n������D��W��zy5��d]	#;�c���P�e��p������rԄ��-��i��}y,^]BEP��l�u�������YC��<����}4�2��}���tW1�Y�C,+���Q��Y��_�{��j���w�~�Ξ9�M�.齆FW�,�X��.�����~�%�O�zWR��L�ڛ�7�5�L��©,��oB�ɗ4B�.8���ڌ��A�iפ���y��(Y�D�פ�arQ�7��G#��E��M9<�tB��2�;��nqCj��"܍�^�!sZ�Vr�7/Z`a�.��rzm���ng>9Z�qp�H�7y)�<��pm[��k�S��=wJ���%�y�wE遇$n��0�L��j�-eK4�,e2c!���\v���t��T��<��D���R᪘�"B:�ع�R��p&�Q�#ykA=ͫ�*������}ϜN��@�� �-XlxV64EB    3864     580��$;`()Ķ�p��&aW)^enc��iX�'yv�e��٨u�C5BC�l��|��Ƃ����[�<��P���H�:xҢ5x��Z��&��5~��{�����L��A\u�9esq�dΟ5;y��,���6��� c�Ǧw��b��	�h���m����!�?̈C�'#ߍ�Mzt�>l��v�=�Љ@���8��1�Ql�	�ZV�W�;R�����ht��'iI�� E;"I�J����r�#�iK��3�$�,+Z�~W.��?-UY�WO�]�hsnl��Ê�X��8��;W�i��Y�!&l�� �������/�D���RUWmF���+��B���!,��ЊZTu@b�X��J#�X�N�����@j�YxF�Z��J��y+����> s��oe�D�7��uE_�y���>)�j+�!��s��4�\�JRS�.�f�1�5� m/+���gy��	o�$�xȭ�L�8*"!��<j��c�
}������#ɼ*�<d����9Vo��������<۷]���^痴�Z�X9 &*�Вh���=�;K9�a�P'��I		�%���z����YgܦDl�p�bM2���r��
*���<Lu3R�;ŷ�?I�,���^��56nFn��BU�5N�p�ٻWAI����!���&�fx���h�g�>�ϙ�w���l��_��A�}�M��Km��#2I9�3i��s�?�C1P���@[���JW\�1h��6��k�����/��3\Z������×Lށ� <A�c�߿�J��q｜�����5D&�=X{߫��E��5o ����W8OH�l	�+v��N#j�}�f�(5���9�I	��ؚr �9�\]v)�~f�*�(N�?̏�R�ɠ��&�{3(�r�?)�����D7R�u���5�F�Ϊ�w�d*vR3(�O�_�*p���	3;��M�lR�$��2���$�\a�4Gn�a�y׌��3o{��'{����/x��bO���@1}p���f�O5,��f�	�E�j�ɣ5G��K)�8P�@!���1?_��c�[N���4�A��r��$ �h��QE�91�jLǰ9���o�f_��LuJ�)����x�A��cGGo��C����#���Cm�?��z����|^������H���I��6���q�ň���⡋F'�h�)�l�ɳ't��S�2���!�$��^�,]�a��K�҆}Go
m��e�z��%.e
\Ƴ
^��9���-�Ʊ���\p"8k�KE���f����ؖdB.���*�ƺ�y�ߋ��۾��O�������;RV���ŜT�Sܥ%�^�-}���L��e��-I�vC�v��R~�����c�=�����	>�{O{����z�5�~肂n���F�Y