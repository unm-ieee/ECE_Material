XlxV64EB    2226     a50��O%��8r;�[Z�^�C��F�d�����c�C�6�"���a�T��@Ψ�Q]�VK��#���:6�YR���!�l���p���vw1i>mcw�.vк=��(��@�tx�ݪ$��~ʊt	�f(�"c��}���?�V�K2�y�<H!�N!�V���܀�2�׽�"�|.qR��YZ���������tG��
7�q��o<�����D����[-.���gj�m�%�b�%SC�h#���02�MA���W���ݕYZ!zo��A��Y�H���	YV/iF`W��]��!�)�Wnrb�=�fÁEGE�T|3-�,hP8�9�#[l�����3`�������b�U?s7�v�M0����w��]0���I�
�;\�C�A��->j� �	V�TIF�����m���6��_AScT��<l~����o�������5��b��>���{炨���x�~F�h�~ʶ�xP=/.˳|�J
����kp�8�w��a�<�3���59�	2G��O#a��wh�Cm,V3���qbޔ�-��éw��B����TG�Ӯأ��.����3ue�؍y,÷�9��b���B��� ��f�̇G����댕��PN�t~tہk}���8�Yp�w��}f	[}�4���k��}s�6Pe�Mȿ�Oi���U
��� A$j3f��O!�?w�y���,A��%*��S�л�k��6�|�MmLp§}��d�N�}`��r񵮫��y��dp~�m��2�zDY��M����z��P��	ʝ���� Aw�Po�����A�S4�?�27�n�	���yC�,\Gn��%p�]-ͩ�ϞqC=�!�M{`�f(�BcE)���Z!E�[s�m;P�4�ƀY��*hjѕ��S�����+��Ø����\��:�d"g�Xa�
����㭖�� �����(Q�}�Onh�S ��<�h蚈�%�2���S�s�A ���|k�r�l��k�!&MH���{�PǨ�d�<��W�J&ھG�m�0n#�
��K_4o��w�9W���Q�s�oc�еvFL ��m�sd�r(��X�<�X^�v�k@F5��ϙ������ap��EA,.��HpO/N<��ګ�]��To�X���"���5���=�q/V\n�!�_qbtL��;N5�I��,�v�7�[�nС�Lq�SxJn���=��C|?D����f�)�.o?�;Z~���̙L9�9ෲ��8GĭPl2���6?�|�֨��]J���.��U\��d�˞?���+��̼Ӣ&�X�s �s�	�	�%7������N�<�wxmz�AS��?����_jDr��[�&����p�KH�)�����m��O�3�*�װʰA��4�}�"��g�:�x�e5�>d�y�ho�����m�GO�#��R�#.��`�H�oX���ɪw�3xVd�9��0�̌�]O�}HMF�t
Sˢ*�%�VnA6i�Gn��A�������aoz��	*
��Й�C`s"Gz�k�KI��L�h�T��,0���܆�6��Pk���c�����ݫ��Y�4�u�-j:%S������ݜ����S���l��(|���u�|0{�q�l~�A��=��=� ,�5�xBpe�rq��ڗ��Ϝ���1#G�g����n��皻ԅ��٘Wx��bq笿au���j���b:�tj�痱 VA[o˵�R�;�� �VG�a���려BK�	��U�LRF�y�������g�
L}.؝�����z����4/�+�Rn�؋�"b�av��"��
�] u�*��6��i";:�_�>��Icʅڬi�g���S=������\}�J��b:��­�6��ө�����ǯOf]���Ld�\�)SJ�ｪ1ÅvN�q�q���a�����k�vo�.?Q����jL��S~_^G�ٻ݆�A�i��5<E�1�Yh�+��������t�#%:3��>��7�ϙ=��q6�iE v��TQ�.�����"Xiv����z��'_�]F�t��T��*��A�p?f��68�ݻw���~�lwപ{�_Ţ��o�LF t R�"J��R��$���X��?:,�@�-�(�������*��c��|wi����v���>�:]����%�VH�h��4@,�P���a�qZ�q�1�xDy�'�%����Rz<9"�
G��xd-u��Liy�3���5 ٹ�T��:$Xat��DYqX/QkH�����"��	@�8�sXj)o"3�G����h��^�{�TR�$�]Z[�\A��I+3;�'��)���쨰oBKC�P�H�����:�1�yxr]�9�2`b������"�U��۬�Z����`�E�Ę2o�;�Ժđ8�o�@z�;*ʝ�Ù=Hފ �b�,D����S��2�1�M����S���΅a�������K�hC����R��:�|�©�`�ʵ�n�g�⇘��'	�+�|�xz �t�>�Y�K��g�*�#��v�
�ɜ��N�4*���nLf*8.�֧�N�e1\+�w� ����RK�<�)F�l��0�niz�m����kW�ӥ��}��