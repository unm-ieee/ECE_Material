XlxV64EB    1c30     a30?�G�)L�6O�om�i�m1��2�[	R��?4:�g�˽= ���3���,�,��c�|͍�M�3�������Ҩ��}��+��|-�0*5�}�K�JZ��"N�'��%��}�]�N�M4�R�O�����۾�x^�p����]�����
!b;٣�� x�vH����rݱ�s��!Y�<!����2kJ8���L�R�m�@!��8�>�^ָ�D��NVo3�QMzj��Jm���L?!T�5�eO>,�Ǻ}d��)��ò�,O{�����{�
���0�	yj�s�A�����1��~3�ɮ�{v{R�ݳ�i�&����>����WE_g��5�p������ퟨ�z�/ꦣx
uV�EF��V�L����w.�N�p�3V�W�c�;5I�SfT�˫!�
Rأ�$~=x/xUaQ����}���������Ҁ�@���sG_7Q�9J�N�z���}�I�������7�w�E�G����ON�k6Q�T-�E�+Z#�y�����pwA�|'A�H˿�=P��6��ܦ��}�Q$��l�BH�jvI�֛e �Ҙ̴�Ϧ�4���SY���h��^n?�\�.�*��+T�f� �W��F D:Y��$�3��C����g��ho�9���{klL9Ц;:��>�g=C��y\x�Yg�5��?��ۖ���X�3�6Lp�V%M>vs��ige1k�h!ߞ��$��]��Z��9W�4���F��;H�6�ip�ɕ@��p�;�J:���a���ɘ�cę���!�+�2r������7/J��f�_k�i�z0��r�4t�b6�l�)i,�?.4Fܪ�:����4�,<����Qm~T�K>�g�[d^^�}����S\ƧLC&~R+--���%���OS�ET�B#����]�c�>�H���Ԝ��0��������
B~�®�oE
�"�����u�HA 2��P|g�?_H��z6?*�k�Ϊ�]y��嫎L���ӇL�9?����!����}}|��	xN�&�f���[c���Ab��p}.	�M�
비S܎J�г]�[<�r�K<!�{��Ȭ�ˊ�]���o����1��Y�z$��O#'Oʲ�VnD���2#C�+W�(摈�8f�I���=��IX���U�б��j{��s��aߩ^�Y{6����Qe[���������Խ�b���HFe��ر�2�B3L��X��j�O�]�,��qט��>V�6L�p��l$s!���I���tTxovMu�,!�<�]봈�8 �uL��2�5> ��{C\�Zza�0��k�pn*�x��I�ad\B!��z~�љ�n��2�N��t���z���;�L� �>"�Fp�O�Ԉ��~����l(ږ �V�&)uv��/L<fVRԙf|�٪����r8h�M��'oЯ�V�dl8�H�!G�;Pvu�� �0�3��`*`/Cɰ�H��"�T|9g�OlRwb���X�lU�K�_��(\��~����*�W� ۇ�{�u��c֍/�XA��	�#��X!��H=	kG.��»����{h����>���W}H���P!���ITҖ��?��9��8���Q�Lͬ|*��!'9
���Wt7�2��D�tMKҤS�}�����ć��|�t�<i$����/�[���Vȱq����f���$�\M����Dݭ���7�y�ģ��@�h�
7���Z��〩;\�p5J^!�m�u6fPt]��立7gL��#�Ր�fd��li�1N�5���&~�I��f��A����?8��T�qL����A��{syxٺ)$#J!\q���_���3���H�=/u�b���s���葇��À���#��S�-f�	W\��N	�w.�.24'����A�I�Z�y�gZ����D˕�5��:p�Iۘ='������9�6�Nm�T{�a��}J�3G▪������I�zhs��5^dKQ�OG �����LB���G8��)TI;����08��S��͙"���D�wC��Lo#������K϶Ǥxn��]ݪeB~��i7�6�t��jO��/�BYu@/������W�$&�H�%�8���Qv�(�KJ����8��Sh�C�&��2x� ��!�������\�D�0�o��B�psd�Y��V�m�t����	7%�먊��C!m�p]��x�,�ؾ?O���ߑ�I�39��F��ҫy����p=ˏZ_daM7~����Y=kҴ�i��,a��_������V����c��1���0�4XK) �.�0*������\"��d�p������Z�b�U<y�e��m �}�JrVs�9�IW\ ���Z-�����(F��#�PJg�ī�	tp*����0r����9l���@!��q�F�(i�y��-��,����.%��2�Y���{K��э�!s�_	����0���e��2u�JW�p��䠭KSڐ1�}9�����[��Co)��$^��6�L�H�t`-s��t��R����I���2���1�oh܄:I�ӑW�t��o��#d�/��:�4!|ays�*7�
�I�YRp��؇"{3.#�����5�&�+��]:Z�u�l[��