XlxV64EB    290d     af0nϲ��a2��y��N��B�Q< 3��j��P����d7~�3`�qMIt},��m��,�{���ԕ��w��n�g���\�uF��j�"�
���쟁R��N�D|;�ڿ��FɌbR�Y:6w"l�����%��m �h��L*�b��^��i:�w]��*F���5�t�0BKs�1���_Z��?��	�Т�^�D.��)A!�F�W�J˞ ��d�|q�5C���E��^���2�������"��� v�Q�M�����q�/��KnW�)�l�å>��s>,`���o���Ktǵ�-+U�ĝ�$d���5�+m�
S���m��H�bκ�BzL7�� *����� ��^�L���F�NВ �O�ߡ�7�����*O⇚9P�k3�@ +�Z�\"/���`�}��J���Pf���g��6���E��|�(�mB���i�Z�T/���M��$uI�@�<|EO�P�ӟ!Pe��3���O�\7.E=�#:D�2B�e#��(�v�_�����1�<����ѓu�E��\�ry�#ɓ03<Qζ3|=�d��R$#)�`ױ��k|�*a�?+!9>�E���o�4[��4E�퀥b�����h8h�#T�$fE��Xzth�^>�������	1�}��:5�J�lxM̓��>���}8����{��f{��x���w�T���x=6s�`D>	SI"���	چ��|��2��u����M�N�t�	":���J4�+u���j��S��*�ġ6���Ԟ5�!�������f���� �h���^����?��M���1��!����`���l��8t@^�(�n�%:G�@&����Ӌ\�}w�G&�&A�uпg�ڑ�Z+��v�4 ��X�x�(��C7�;|��p��JG���3�{��� N�oH��G�ɗ���t������4�qO?7�^� �U���=,��j�ۄ#��~@QnR�l��GS�M���Y=5y,J	�"����>;RT~��z�gi�?�j>��գ�L��)�~���y�P�ޠ֧���zCz�`T^�WZ����`8+�r	�$d��6Z��p���L5���r�v�dOY��N�>�8��܀Q����g�������y�����~o�	S:I\K|&�wc1ρ�t��be�{ʺ�����̈́i'�M}]�>3�ȓ1�T}���Y�N�3v�{Q���<ͼ�Ga\���R����|8>M`�V}������m?�4A�C�L��ا5��}P^W1�.V������������}��
��!�oh^P�;;�g�:^;y8)��=��/]���+ �?Y���c�S+�*hq<Ơ*�z�������s.����0N����S���w���c�F�R���,�렞�Ų}�<7<���	�HSoE�H9Q:8M5a���b�҆2!ο�=��r����[W��a�P��Z��]�)%�0z�}x�S�I{���$7|OT(�FU�a76�x�5l9h�tj����'B0��C4��ƈ��º�'����܇ILz�Kd~��S,4x��f������)i�q��n.�틠��ʂ�qu2ZF��������]/��϶�x�`�G�+��l��kW�Z-��\+|���UP��*�a�� ��È]"�Vk��s�F�0�u�t�
�1�-!�,f/QP�0���X��Đ��"I5�45L������]�g�h���.o<4� �^|���Πk�F�7Lbut1R\����w��*!P����=��K�*K��B�\ډ�K��Vp��\�KX)�0	��_Y�9��VP1�D쉃J@`�eFgڗf��/����q'8�=?�?� P�oǶn�R'((ko[QwE��
f��PT���������*�s�-.��m�4<3�7��5�3#q���U�fe5�(�dL�(�ӆ�7U?�x��=1�ڰz���g{X���XI�x�dN����!�=a:��n�f>Z�U��7��x�H���N����
��S`~u�FxC��|}�2��yk3#�:��<N��H��͓��vݱt��+i���)C�8�#�t f�}��'�b�L'+��Y�	��Q�g�W��#aV��L*6O�J�xR���o*�b?�"R���CGcf��!{��-��x��}!L,+&DʾA�W�<K3��{�J�v���cWlu;$L��3�G��҄���^�����WY` L���fw�u����Y/�]����+�`@.9�ɠ���F�x�DWfEu�g+C�dw���p�IUX
�'2	4�R�ε�y�PI%�[&�ǵ�PD�|�����F���k6Yi��\d'99%)��d��mU�A�m�bXu�Hy�^�Esm2��9�"���|��4Я���N�M�v��&����2v��yc�H=�7��ѓI�*�I�*����?��P��\<H�GJkܥ+��U�$�	�֕��2�����q�h����_��D.O$�Ѡ��Q�m�pKbZ�6V`)�]㺱�#�0⌹l֟ �%�$�?f��T���c�L�l8�f�� Q,Bɷ<��N�����۶���Ъ�sD9�u ���EȠ��!7��or��d��;mѤ\x�pl՛9��ta23cp8\�x�'9�� �än�w.z&֣�\�d�=��@���HΜ��Er�Ӈ�_/�Wu�� J�j�emD��1��h�a����3���~���HE�>��Z俴�T�髳��� #�n�Uy��gi2z�<�#H�>�A���������9�_ͭ�x�P�I|��)Q"FE�rN�AV�m�r�@��x