entation="horizontal" >0</ScrollbarPosition>
      <ViewHeaderState orientation="horizontal" >000000ff00000000000000010000000100000000000000000000000000000000020200000001000000010000006400000141000000020000000000000000000000000200000064ffffffff000000810000000300000002000001410000000100000003000000000000000100000003</ViewHeaderState>
      <UserChangedColumnWidths orientation="horizontal" >true</UserChangedColumnWidths>
      <CurrentItem>ATB_MIPS_ALU - ATB_MIPS_ALU (E:/ECE.CLASSES/ECE438/FirstHomework/atb_ALU.vhd)</CurrentItem>
   </ItemView>
   <ItemView engineview="BehavioralSim" sourcetype="" guiview="Process" >
      <ClosedNodes>
         <ClosedNodesVersion>1</ClosedNodesVersion>
         <ClosedNode>Design Utilities/Compile HDL Simulation Libraries</ClosedNode>
      </ClosedNodes>
      <SelectedItems>
         <SelectedItem>Design Utilities</SelectedItem>
      </SelectedItems>
      <ScrollbarPosition orientation="vertical" >0</ScrollbarPosition>
      <ScrollbarPosition orientation="horizontal" >0</ScrollbarPosition>
      <ViewHeaderState orientation="horizontal" >000000ff000000000000000100000001000000000000000000000000000000000000000000000000f6000000010000000100000000000000000000000064ffffffff000000810000000000000001000000f60000000100000000</ViewHeaderState>
      <UserChangedColumnWidths orientation="horizontal" >false</UserChangedColumnWidths>
      <CurrentItem>Design Utilities</CurrentItem>
   </ItemView>
   <ItemView engineview="BehavioralSim" sourcetype="DESUT_VHDL_ARCHITECTURE" guiview="Process" >
      <ClosedNodes>
         <ClosedNodesVersion>1</ClosedNodesVersion>
      </ClosedNodes>
      <SelectedItems>
         <SelectedItem></SelectedItem>
      </SelectedItems>
      <ScrollbarPosition orientation="vertical" >0</ScrollbarPosition>
      <ScrollbarPosition orientation="horizontal" >0</ScrollbarPosition>
      <ViewHeaderState orientation="horizontal" >000000ff000000000000000100000001000000000000000000000000000000000000000000000000f6000000010000000100000000000000000000000064ffffffff000000810000000000000001000000f60000000100000000</ViewHeaderState>
      <UserChangedColumnWidths orientation="horizontal" >false</UserChangedColumnWidths>
      <CurrentItem></CurrentItem>
   </ItemView>
   <SourceProcessView>000000ff000000000000000200000159000000eb01000000040100000002</SourceProcessView>
   <CurrentView>Behavioral Simulation</CurrentView>
   <ItemView engineview="SynthesisOnly" sourcetype="DESUT_VHDL_ARCHITECTURE" guiview="Process" >
      <ClosedNodes>
         <ClosedNodesVersion>1</ClosedNodesVersion>
         <ClosedNode>Configure Target Device</ClosedNode>
         <ClosedNode>Implement Design/Map/Generate Post-Map Static Timing</ClosedNode>
         <ClosedNode>Implement Design/Place &amp; Route/Back-annotate Pin Locations</ClosedNode>
         <ClosedNode>Implement Design/Place &amp; Route/Generate IBIS Model</ClosedNode>
         <ClosedNode>Implement Design/Place &amp; Route/Generate Post-Place &amp; Route Static Timing</ClosedNode>
      </ClosedNodes>
      <SelectedItems>
         <SelectedItem></SelectedItem>
      </SelectedItems>
      <ScrollbarPosition orientation="vertical" >0</ScrollbarPosition>
      <ScrollbarPosition orientation="horizontal" >0</ScrollbarPosition>
      <ViewHeaderState orientation="horizontal" >000000ff000000000000000100000001000000000000000000000000000000000000000000000000e6000000010000000100000000000000000000000064ffffffff000000810000000000000001000000e60000000100000000</ViewHeaderState>
      <UserChangedColumnWidths orienta