XlxV64EB    fa00    2cf07B3��$꽜���@����X�@o+͎�fYo1K
�^�)I� r��2X��>�܏="��w^��4�t\��ݢ}��Z:�Oi��^E �/����-���\1�\F����3����?EX�W!kG��Y)b�{^Av{v��q�'��[۰L,�u�J�Y�4HA�{<�k�����1M�iZ�H!�J����~�������/Tr���s���L�cm�Je��T�{
�c��3�H�+�j
4�i}���8�j[kڈ�c���=�5G�n15�w���;�1�E��2B�m"Ph����Es�r�ʖ��ww�F�@T����g�<���`�y���˸�V|�b'�Y��{��H�O(�8��)�
�n)ͣUfN���g�Ug����?���ќ~����GJ:d���Ip�e�%Z����h"Z�߳�ϟ���E�>�#k�Ժ��S���7���� c44�)a���Q��QP�]�����Nĩ�h2�؅G�43ޟ�1�R[�,�R��U9�n�9��z_~��A��Xpf��G�㇠^�(�&|�O��$b1�Ƶ
���t2]ܩ@oR�C���2���@���z�W�U��_��0��H���Bv<�f7�B��c��e���V��_�ta�|��(d���A�61k�j��>�!�Ɯ�2!�"U�^+�$f�7�V�r�>.+�g������]���ns�k>���/��ލ��U��W���j|c�Ҷ���{�.�� �*���~�1+���T!�L���->�rgT,����F�՚7��.���>�v�d3��8�D�(v ^�:h�
�	�b��@.�2Y�<B�$��ƈ̀ڿ�ٯ�R+c�,ç����X�;�P������}�/��K>rJ��%@�W�ż��ngn���� ���~(fT��i|��E�	�9��"�I��fRf����k���J��5�>c��T"�'��{i���"<Bݓ��gJ�䱊��C��^����_������Φ�w�x��V��8�����'�;s�5��5y�S��]Wmn���\��<�lB��?�D?��GA�'ю'�+'��$I���)���4���L۠��%����62ø�H9�θ?g�@�D˴�E���H�$(R���6�ч���GK�G#P��۪�5���4.���4�'�O�#��I�-�u-�RNs�u���W{|�6L�lFy���zӚsXGl6mI(���X����h��Ae�V(�q��2�5c��P��&yӁ5�rӵ�mT~ m�@V�g7��?#�ɑ���5Y!u�s�BN2U4G,��*s�B}�*�Cctr�"�{%^��(�]Gg�(�7�`e���5���	kL6���X�:��X�%�4�s�����`�]��n�[�6����8�F2��ʝՑjxp�x�&E��[��-�~��=�uH�v`n(��cT ��(�����'�� f����.�^r�N�:��u�X��^�HB!�����Da�H��?����8��\��G����<6�mr$�W�Ǝ�Vw��ʣ�6u���%�j��jY�z��|[�����+O��;����#�HqsM�*�-U�K�*X����L�;�=@�Ѯ�ϵf�s�w�_?�9�$���+������!�5����_?�%�X1�
�Q��$:.��W}X�`Q�U����s�n�xYT�X������ܳ�Q�xc���s�:��^��~��I�oe+�̟�=���0n#5G�M}u#K2��ܐ؟ŝsT|jn����F�\�w�h������!iw6�^����SvG%����Db;00�c�䉱��)W5�,�3�"�G�Ԟ)��E���&ng��0�4����?�P�Z�����7�Z� ��Vo	M�}u^yX����ϊ�|~��\�!�<Ӆ��	W��έS&�b6X(�F��	�4�.[%co�i�/�c����C�z�/3��D�����,�Wø枕زϨ�� �+��I\q��X��D&�-. �>��N�&��a��[ev��44�����x�lއmK�x�y��[�r��R����]�XfH+/�ǎK�v9q7�^ެe�?��%�T��z��7�䅺�\gz��f=�H���^��|\F@�R��[���7�}����U��U�����Ƌ~�!��	ce�z��l1��vs������h�
��P`�N�==��Nd8:>����4�"*��	.h��ҥ��)�����<�2oY��kjϥ�<��C�f!9�ِy?�{�l{��!�p�Ӯރ�pM$����aOQ���x5�S���ej�<u�e�g�����e�*����R��A��շa��;���rk��>���rP�\�x9��kQ'�"}�!Wk�!8ܔ��P��|����#yjlu�ċM�+|衈2����hy�'T� ,�A�v%8�L�JW&@�7r������M���S7&1�����)�����!�bM,����0�yS��"4vc+���Dk	yv��)��<񪖥��%��N p�<�yB�ۀD��h���pR$�����wf�QxmECU9��+?�jJ��wS�f6c����.���Z�C�h�Iy�L=���=�����}4㻗�Sʐ��h�>�k�!e��en-:M��ɂ�XI��1m���I�
�����3=ޙ��T�§f ~����ƾ- |fC���g��[�vx�)T,zF�jvJ�#R��8��K� l��/�bp~�q���SL&o��w+�X��72�Nu9	�F���`	���B4��!��7���î�T#S|H���Z��V���z��ߦJ`|������R��/�;��g���m�����L�#��o �ܶ�	���T�=�pt.{R�aC�B
�������jA��V�+�A>�?��h �`?<�~4�G�V���^1~ukv�������ږ��̪�sC��W�:�h���ּ�*IL����;��q.����PL<�=xDO6��4?@��=���_�S���E g"�}�u��j��ѵ���׷%���l�;�r�iTH&���3�}�#{��^N�Z�-�B*AD�;!uL�3��K�Fi^�����h�W�G'��n����/{��&*F�{1;�)�4��f�=�(o,��bp0�H:���(�9�>DS�3��X#ֳ��/=5��69�5$���D-�r{jd!f�?�ǖ5���ΏՏa�t��W� 1�qӃ�ak�k��,���i���1��5��;v��C%C�~:L����
O�c}
;'֣����
�6R��`ֿ ������ԉrX���ɮ��b�-��(�^7�LGa����}�3Òl�p�y?��ހB�!a�k�e|������hz?�DD�EJf"~�����;sݧ�aOǂ�H���hI�h���R˦�35i�{�&�0�-s8ڙ���UJ�((Uؗ�H�^b��V$�fŁ~�Nt��6҈�Bs�FFv�������	�ª5��-��XX�z-��}�z��g�����b�����j�o_���-EU��*�Ũ�+JO�mo`9B���ׅ�E��8����Eu_�o�'�CG� a)�Cvt���ט�Y���
�q��5J�,N;������F�6j�.��c��ny3�¿s$b����H��
d����?\fm�%0�4`4��+$:�3���̯~7��xp�?�7�|��^|><�LݯSaK��������ɢf�g�%�K�������lZ��@bg�M�����0��u�͞�ՋZ��!��tW�J�CCҟ�ōe�>�U��V�2=Z&��
��!������Q���H(" �2��N��	lzl.��hA��ZC�k�O�NMޙ����h,I��^:����S���L�YR5q�`7z(��c��)e��耻�DXӂa���OV�	��=Ɗ�2s*O���^Ѡ�6�;����� g���7-'�-����T��L�y�?JA!``=��a�S�:>L~�5��Y�u���_?�o�̵8o�5H�M�>n�U�֍�@"���8������[n�˵���D[x3�>@�9�CB�M���ܽqV���۶��`?X]{�Hi�ث%��4���н��$+��/JdII�� @W2�x�S�:�sRQ���.O'��e��&�-6$~���± ��ysu���=��h�ay?FK�kZ3}]�	�s,�p7��(Y�Z��� #g�/gb@`�߁OXe�3�o���/���Z�^�l�>�izuM����HE��&�vQ��Y��H�,�Fɧ�~L��(_�ĕ���e
ْ��0(����MN��F~'���7��$t�9e���E��&�w#�2,�Y����$��q�<���`��Ad�]a���m!i� ~��2��j�9��-��؛0(՚N���%�X.�*�{�����$�>ѧ��A�}r�+]�ᓇT���~��u�X�3*UG��)�@�R�神|G�%�^�����x�)_J�� l�WϷl�>���qH��F4�g�ZBjH�K�˅�m"��Յ�,�h6I�|�=qb?���z.�{���e��~M@4Kz�8@����#@+MK�h�$�Y�"-�u+ ��SfPk\��`��&'r)dn�ר���]:5+��V����=�)�V+{kt�Q�9�4@����9l��rpU?S4UN��T�<��fR�y�Z��B/WS���ԇO�|n���}A�"6�-�&;&G`\����b�[/R�t�D�&�:���(�Kf�э�TX-עC�n��`-Ҍ�a��'VH��f� tV,��k�4{�c�oF��<�d�W�qJ��Z�5'�'�Y����߾�E)�RbJ���c�|Z�.*2�N�ZQv��� 3H0>�����{��~y�j(h쥙�7x;�&x��$='p�S
y���ߙp��՛�2�&���������9��maB �թu�]x'��?a�s�-��l�!
*���kD���	ش��A�e�q2��"�(X�q}�՟�)�2B��"bx�&h�qs���_�
H9F! Aإ����;<�^G�����|9�Vir���������/+�*y�j���YY�oI���z
��X7������݌��Us�ۚJ��jK�Ά�Osq�P0��.�L���O�_��S+a���P{����.����tc�x3��^��~�Cw�V����ԝ�'���R{ߝD7��JJ�$�6#߀�ٔ�?5���_��S��dg��V�F�_�u5?k90<�s�H�r�	rm���Ew�:�n\�'�ӱ�#�0-�4���Q�x�f���z�_���Y��N!@!s���I!��*VX�����~2����L�c����܍����J
�&r�Y�&�a�1w����p�o����T�f�!<�;lyu=��F�;��ƾ��O���������u��hz���]!N=U���;x��,� ���tr/;�n
-�DUM�_��e�%;]96:�Zפ,��ԁ��莭�E��2�����r*+���o�����HƺZصv*-����&U�<sJtPl����3������:�&/&v
�﮿"�J�m`K�Yv�^�V��\�zJˍ���Zf�Nѷh���?=�?[��#e��d�a�1��Dr�鬺��-�\)�j� E����.��60n�2�J�ɨ��_ޏ+��h5���l�uzM	ǣ�oXw���E����Q�"Ć�OHEN�h>�K�K`	#R��ò�q~���'��PϚ���+��θo��!��"���kR�}��~;��/�}��`�5F'�EZ;%a�U���R���b��"���7���c�TjB�c�(*b��Aݵ�i��%>	16�"��o�m�'AZ)�E����q�Vɼ�Z;���K��D᝟���gS�w{�1&B���z�S�ػ�f�@>�ʸ���V�4��G���4���������FʝUL�J9-�!�t6��W�2|���7��/�ӻ�����	E,\A�5U%����PCSټ�L��b� �Ȋ�\�!'�/T�IkP�������C@{� k6}�^g�[D�[@�4�a��/���n�[!+Wn��8��@���)|�����lV�!���)�C�)��d=�^��V��>�*�vF=��j��Q�M�p[�fg8�w<�����1N��Qw�)�"�XZ�LC�c�|���wyk�Y�S����i��X�h�x���Q����������A���$�j����	���lT+����$�����af��ʠ�]�;�:`v�����!f�D���R�]S�n�Z�W(����oS4֕������<��J�'-o�����.�J(�C�������@���r#�jڂ��!6���y|Ê��������:�G/��$���1��ws 9��Y��E�X<���/��~�A�օ�}K���,|��{�sr��	�M���Y�t_��;��݁dNr�f�틜�-l:��n�ճ���M����`�2��h��بeU������qYW�Y��*ڀ�댼�2�����|�a)QIy�S�b��n㬛���A^�[��KP՝V��x�B�3�S�8L\b�|�^$��ل��n�L\�'��H؞�SW9�.�������� ;	g��b(�ˀQ�D��E�sߚMk����VT�4�1�0�8��"�a,pYg2�mz��]��������n��핚S�#�>�/ף$�ǰ�3����:F��e���Љ�pz8��-�ֱ_6��B���<2�Nm�`���p��8���A��-¹s�>YKO4����_lP��>�8�L�6��p@�����y���0�2ih=��꧆u�:D�vO�~Y��a�@��R`?CA�"���<F�P�s���Kv�3�Ѐ�EC:>-Tሢ?@���bBm�U{�&Vիd���H�-��mK�@+{�=B�Q&�Ʊ�sX`��A� zI���"��@�!����?~ �;DW��>��N�JlF��r�P�ݭ�>Z�SV7i�-�R����,����:�����ox-�W�ʌ��IlǸ'�]ɹ�C���"�A�ǐ��������l?����!a��X,q�YcQԥLߌ��T�!�a��}c5�*�Mg��/����H����/����B���1���`b�^�ts����������cPI�1�+o��6oO=rP���ӗ���$�)�aQ�O!���Yx\�E�G!Mh9�L@��Ɍw{B?XВj��"�˿1���A�x؞*T�;�v��(l�݇_ե��mp1v��P(M*�D�ƅ�.@+�+%.
�I;���Qv ���ߌ��m�3�L8r��ݸĭ�&�}l=#�����:�dZ��3�p-R��	a��+N��n�X��>cb��(pe�d��\��ԗ���:|�vE!��Ό�$�3I�FM�}:�(]5F�#�{����cܹ��:և��Ë��=�F5��Vzα˖�As�"{y��	��vE��!�����$0"�ZUvG��s.�F������-����s��t�]�nL�Ν���4�B��w����9>�Ê�g>E>I!Y��^KF`ӧ^7s�W�(s}�&���F=$�H�n�EJ�9p-��4נ�0:�İ5�?�2�<����~���^$٨	�	'csg�F0��=T��)U���aS�IFVÎ�Q+�֙��H����X��|��ņ��'�8���5�;�"���� 
Л:,&��Å�#"�P[}xቻ9�M��V�1��YA���B�l� ile�&������9�{7��c^��ꊉ��$�� #4@�eH�	����tqI,`�p�{��J�O���y�����w%j�n��I[�T8�Yr���d�Y	s7�q��)}:��`M-�����τ�
^��UXچ�5�i���u��۶�m;��l�e�N'!���f�UE��R�f#Z�|��6�Fd�h�S��=������:�+���.�	�x6�\��H����Zp��"ZǠV��L�������j=	�c��Z��a~V�Y��T\z�K4Z\(�(; � 9�=�g��P�2���4�tìG�@~Um{����T������z�$��7�k���H�+�fҦ?]B@�׫����*5!�#CT�A�������Vqc�G�2'����o
����KD�׬��]nj+{:=yM��.{;$gݵ��,M�3�%&h�ٓ���ꊍ��U��0��@3ۘN�h�����#C��E��G��&�Fܜ�Z,�^t�~	�^����T� G���ИR*�$��ϫIӎ���`��w���Q�o)���D���Z�-rq���I��!ڥ.ş+c2t6�Mi)����,�w�fa$�\��s7�����i:oe/?���M�7�7���]ͫ _�u'sz�����X�c��cq'�[����8�5s���|����q�(q�W�v���aس������X6;�	[i���sb�����s`Urj�PR��[3e�-������̙CM=�43M�~{����S��޲�ڮ�S���%��8D��_�3�?'����_t�10�l;=�[g����7��������U�*��r��f�e�
\�������W�J�~H�v�sdM���F\S�}1���=���Yv�/��{�4E���"���_������q�9!p�>ʿv���ӑ���R�a�崸� #_E�p֘Th��������}�F}	���Re��|@�0\ 6��t�I�c��a-)]>�/��L��ށU4�/���\?1C�ڇ;P�<}oS(c&����cz�V��wۃ��x}��xz��$�S�t��d�S9M�>��Cb��	�MtG��/�@Hv��-�|z�@����&7�E���]�HG�,R�l�1}�$[�m�E���'gd�<5&�
��$>�
̪F�7|��N�8��qb矷-���������t_�,�Y�#�긔�̲2;�H)<}�/z%���ZJ�Ppi\s.F�5�.��7q�
�	Ff����#)��#�,��j��ظ��Jٷ7��&�&�a{l\:���k�U��6�������'�}�Y_X��h��4(<�K�������M�	�21BC��- 貉wkRx�
#��1�>* b*^
����4��e�,�6��ٵ������?�	tcE�7��e^��C��k?�7X�vw�X�sqv8E24X����sQ��A������"�f@���b��?ͻYk�'��Uw��tc���*/��5u�"j �2��a�O�\����5��/�󊦆ͽ�C�$]��;��E���N{�_K x^Z��I����f��t~�C�**� �|5�E�z:��~(z;�ʂP4�}3A�h�L^���&{!i�e���7)� �G�ܤwA:H����nTE�{��2�>�ePjڜr��=�J����6���Y��`/�%.����&���h��$r�_rpa~�K�y�0q0������ ����]!F�����͐f���CJ8�ouچ\��lQ��0�o���K�K�2�����M����ԅ�����P'a�����j���AS��2(<����\��"�@E�^+�y벹Z<C���7�^�)(h��Zq������Q��V+�G��ȦOw�Ox]8+'�m$vx���AH2V�q�7���|�C���`���9�A ��CA||���r�Qti�2?NH��ⓙ3�f���R`:t� "��<Η�HA��֏&4�n���@v ԗJ7'ԆbĖ˨����D���Q��c���L����!f֚����y,Vc,{*�!�㚧´c�E`s﹔n5��a�~<��������J'�$�?�)zŕ��sFC�_ړ9w���{�������`ށ��B�������tP��#�R�����-5i�����9���Y�߫|�!l֖U)���9H,:�)�.oʍC���u���jA�^!����p���rp�Ĥü3o�W�������Z�a�oΑvv�"��E���#0�p0#�Eg�{m?@�/���Y��7׭VX��d�����qn�Ev�*G˗��*����Kb�O���. �b�����W��P�^KԵ�4Dc�ڿ��e5"�F��?��	�Kc��e��L��_���"�~��h=	��p������AP��BM6[[i�L\�ʁ�7���H�(��p���8�,����8	��\�����Z �;�t��nY�J�YH�Kc��1,Qx�<�Ҕ�J�-����GuC/�3m�{�m�[�������	QS[%c�wqC������l��
Ԭ���,X7[�΋��;�w����B�4=��r�9�6[v���+\�> h��}o_<|�)��+�HO��#q$ǥ6�,�56���q,�<���6+�N����1 ��x��*�}�o�SGS�3�z��ͷ�Ê>���z�G7B]/�q�b���O����J�<	������r7D��ő2��	_wX_�h���Z�֛��='�bA~��:#x��j�Lm<d��3���3b�X3�q�,���,��wA���i+K�C�@3�p(ha5���ķ�P��]f��Z�/g�����E���)�$L���k���&5�->O(Q)1�i(��v��az����d҂�
v���w��C�ގꜫ�ĐO�SY�(��(��Ml�
�sy�WX�]�^nf����_����QVYO��B�=A]bt%a?uy'�����ƽ0�y$�H��%}�0�O#=��a���e�|1�Й�	�:eY"F����)��Y��foa�d�_�(��0�/*��vF�=JʕL���G5[��;d{�^c��a�+�i�}�n�p6.H��5Gx��.�>�VN���N����.M��)F(���2o�U�G�
`�DR���� g���I��g�����<J2���_Bb��Cq�A�j<��PD��������$�b8�ˎ�{�)Z��)s �����U����"n����5K�8ZF홣BEZ*�c����C�r��k�S�z��۫�M��Lf�k�P� `���Q�Kᜋ���D�
5��XsT��-�����Ԇj��)��^R�/r6-fV|�	�?A3�f>Wona�.�$��C9��;�D�����`K�;lQ^MYF�6&X�aXY��J�3N@]q0u���8��v�RޜϰT����0HF� &&{����,���x��y�x�]�Lm�K�'��rL�{�-�~o2�KN�
�j���A��47�"j���:7#�Z�nI����%T���6+�¼3y���hX`�5!x��<#]	=���9s�� c#�ى'��5�?�s��y ���J�XlxV64EB    c805    1710H��\��S�-|���f�8j��)e`M��2���-�PI}B�qF�!Bρ;W}l��Vx�Ʒi�\��/!m�(�WC�3�]�E�J&p�}��{N"��Q��~o�iJ�m�/���.P��0سZI�L�kBe2z!\�Nt��yV�����X����^ψ���/7f��{��v^�ׅ`y����GH��R��#�Ʈ��:�-(\WH�j����)t�(y[V�C�25(C{��\-��1�JX���؇p��~Vr��h��jN=U7{;�����g���G���[���;YH̲�����(�����B��i+�*�5��0D5�����Ԥ�y��:b4;�Y>.W��@���5�"�l�R�|���meI���?���N��_����c���]��0��m�Ȍ������aݻ�Q�/'��1E�\�c2�������q�Uʙ�Ic�Y�,߉ԍ��0�֩-�g�(|�)<�+hLf���c��X� �$y����J���!�-g��}�V�����WO}y�1��	����]�<�
h�%���tv =O{!�U�~ֽ��>;K.������b��_?�yR�>�kXbU�L�J��{P5	X*3��v耴��B�̓9F���{&��X�C�l`$��`O3۝�<�hܲa���'vgL�V��b��[�Z)Q��_�>D��|�]SX�k}�U/uq�����R!�J�9��/��|2a��I�����=Z��!��>'c�[&OU�*��#���-������Or����5�j��|6R��t��W30�<�8�kΨI�[��-�v�--m�>��B�+�~4�z6(�@%���(^Ad�rO�k�+��G�pA��s&" �?mj"ƶ���z�A"��Wc�[��X�~/].$m�1Ȗ�u��Ό4~`rq �	B��[ը�A�nx����2�7@�;%���v8�W���c 	����Ľ6»���i9�����t�|ŦOq�c1�?z�C�5��
U���BĦ��8l��&�H�q�?;g�䋓~Qiz�#�:Ed�"�A)v�،>Cط?}�<����b�D�IwVzh�P<���� w�l����!��,t�c���j�[��H[�L�(��F�p����LM��M�A� ����Q���`ɧN:������|���G7����x��߇3�>�;�`�b!!V�]��7�^&W33������Q¬rZ<kM��Q'3��+���n� O��9�m�O�a��Ғ�Dz(�k�J��u/����o,�y�G� .3iD(���\��5��q@=f�������W�{����-���WZQ�R�ܸ��-�q��KN.�7��7
�ik����h��@����6Hi�R%�����-����y�d*�Hn����o����d
.���:�.���Y���y�6!F���A�Xi(�#a��Mr�2��e����{c��w��nϸ�_)�����
[2:쎑_��N�w�H�=���m����������%\1h�7/7�x��j�|�!}�%Ŋ�wYv�^#�}W�}Y$=�B�4cK:O���j�C ��ơ&�-l<�j��랽8�B��v̰S��o	:#�;))ҟ��$��3O*��#����H@�ZH�(��cp�𛔻�	ˬ���xy���C��WXFȵ�ϵ�Č;a ?���B �S�%�¾c�Zh�	U�cl	������rr�Z��R��&U��u	yd)��Wx5�
��p���[�lV�zT:K~�\��t2	���\`���>ō8TM�k�~�(�V���?x���8
T٭5�򀥴���m�o�^X�2�q|0����� ���1,bV�&݄�h�zl���[~bÄ �m����כ,�>��(�2iL�e�A��6�.1Qj �ꂽ`J+����p`;��$�6ut����O�:�q�>&��2{��Q��n?Z}�r'�~ܽ��~�~��iR�6Z��-�bk�i�=��3��堋��ˆ�{3;�kU��Ů���ʰFU�a�h�*��\b1^fb�J�]f�4*��f��MǕ���:ϗ`#�*��8��'����VIQ^`O�[���WͯG��
��QvH���A��e�ubu���;T䁉ͮ).LJ��VE216��>=�L��V3����i���z�^��^:/0�:%�}��T����K_�VM-R%�q��be�V�e>��?�ݪ+�ؑ ����d��P�=-�9��Nñm4Q����,�f�F���>�}q���d���?eJ�U��Έ">� Ro@����]�}��>��f_�l�'W��S^�����&eբ*���)\�К��\��U�1��x�B㮬�!��*�ϫ��Ň.���s��
��qE���΅~��]�n 1C�.��XieM�SW�f�{�J�A0z��)���8���@�9�Z�	�?���,�L�ȕ��8��.U��.�?�m�4H}��.�kX�@�TS����T�����F���!���x-�-BGt��a��s�'/@�a�ߩ�"HK�hF9
v��-FӰ#EJo0q��A��J���"�jC��_jܫ�^(� ��ۯ�B�J|���M3�
�&�7^��q9!%Р�n��bm��#Q��t�7�����pU��ʚ	��R�S����5�7��r7��bk�>�d˒��̎!�x�%e�_friyHG�\L��W�v]��y1e�8VJIV��HG�'c���I��[�Bd�������D�<<%k�w�Xg��d�T��Q�g3mH��!�~f�]�����n)`ί0��(��S��fC�~���n�7��6T�'	���3pa���p8��s���{�?�U	0�J�t��~�'bv:
�0�\����^0Cl:Nq#k�ʦ[K �8��JOR�cL����p6�^R'�O��ȬM��6I�2q�����N�ݼ����
\��<N��h���y� �ٚ�H���0ؿ&_�o��/1#茔M#�J��A�d��cu;���t#u㬡�%���-=t�G{����´�;*o^b>�8�.��~�u2����.Y��(��Ն3h�Z�l�����T60	yjRہ��)��O{�f ��H02����I_�0� �|��~tŹC_�}ҖL�=%^zط�V)"�c�T��9���d�R���T������څ��g��>I97���['�>T�#l��En���;�6Ҿ� }^�:*�&Y�׬ӟb��+`F ���|j�N�Ī���72^۳�$�HC��4�����k�����h�*a��C��������U{���G4� �Ƃa��� �Qwq2�=���y"?�*mgՆ����G3I�u^�-��<:��pbӤ4i�����4�>���^q&�5�4��8G��v(O���	En+��K�����̝���T���/փ���8s�`��K��
��9b8��?���6��Jm�P�=�  �.;�L�e��ɽic��}>��y�i3�|K�_�Û_{�qxB?h�5^w�?+��@m�:g;�D�Q:���"�������1���rqYp�Ř��B�b������ZP������}9HC�yH	>5]�8�2(.?w"$��j.����в�4���b�a���q�H�+#<,��<�n���5!S��S�,>����k�Ե�'��� �����m��1���8¬�n�d�� 4�0T��mY�-B���xh�]~5�m�qj�'{����@Jk0�m{����Q	��mZ�����W�5�o���lWg��b��k���e����2��ߩ0X�h���^�;U��)��< P�e�۟�_��Tɋ܍?�0�#~X����V�hW!����΢�ﾺ�s>��%'G�n_�&����p~�^�|8Z�Ђcۢ�;��	���*��������ݏ-��bB
&�i���#�ekY�d`S�0���o��E~ �A&��E�L��U@<��6ڥ���?��&���|&�����Tvo�p:�&�o�JDGn��a
e�xu�e����n.mbPf�֑R>z�EY�D�~˾���VQ��3����[�z㽀3u�?��W��/Ӆ���I��o ���tf�Yq�[ZS ��������͝�,�
VD���c�IY�̤����V���tclp�aa(K���a�R�6�H���K�&�$Y?�l�G9�� ��a�j��՛�9'	�ȝ��F�$\Ue71��Ҍ�]��V���j��;�s>淇�3���`p�tHp�,~�;9��G���A�!�`_)OW@�i�U㷌�(�t����Yᕠ������e�-�O�Z���V���f�{aCa�=A=�_�	�/	�B�2+/��?��6���mˡX��P��4�Lw�X�lqՏIJk��,P
���Y�����S��T�J	�<�e@n-9^�bN���0;��EH�W�6���`~臕�t��/�K��c� �����w���6ڑ^�k�U2}u�'����FN�uX7��k�wf�$d��E�9�� H�?S����m��,S��ֲj���y����r]FQ��<^B��0 �	%��Fȡ��.y˙�dc_�-Z_�W@eC����*�n��s0-�t/�I.�Ho[�>�z������?C/]o�o�ů��̷������~Ք� ���}� �>rNa���쩏*Sh��ӐĠ~{���gJto-��βHBI��e�[Kҙ�_��MŮ����L\�p�x�M�������V3H�$� ���u�S��1���0s]�z!PŎ�u�E�2�@�`$�
���,��E�#>kezQ�GIkC��=��w9Ч1:�/�/ߛD0�m�Z���>[/�G��i�Pa��ގ�͏�%:SP����� Ы��u�NAb�(U~H��#��Lq=a���(z��H�|��4ҏ��������#v�Aw�(c+tW&:���+����P��b�Mg˖�?,Z��u;h��Yt�wѧ�r�.��P@�D�6�F�+��W���q�/d���`��ZdD,�}J��B��$Ơ�W/���ɗ��d[j��dkc�C�**v�/���,�B���R�f�-�@A���h��,�����p�9s���
�<{�������������_�a��Y_��>�r01�j d��hh�
4Q��!�ivKw��	�f�~��,�0o���̎�����Z��$�v���a�\��Y�%�JNx��ԩpu1�Y(�i�G({�R u�;�"`�39e�oIk
=�4ɦD�<<�"�� ��i��B�)5jx~u�(H���Q�L�ko]K��[���B'>f3�{�{����I�GLQ>ŸU�,��v���UI���PB����Ⱦ�Q�k�^�O�d&�]5�=�g�� ����Doq��ע�"��c��� 8�c�T����%6'�9�I
�W�d���w�&I��6��ӌe��;��4�Vl�����\q3���
��O l��9���j���.��Ux�j1�h�r�Ȇ? @޾;�����6�}F��@�h�)�m�H*ZT��ܿ�&�O����\�H�@�͎ �]�2=�5�Y1�o��՚�zs7�@$�e�Q��<�gy�P��sk���QI�?C����E�3AKT1�Q��1#��b��{2��n��ŗ��"\L�N�6-5�8 �ٸF�@��A�M�-.��(\n�}��ٻ_�)<�\��0�!fK�m��l#��I��j��k+=��uK!�J�x��h�nW���؝�>�M�lL�5K�GA���7f,��֝~����6byt6�."9�l���²A������Aﱶ��{�