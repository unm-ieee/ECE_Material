

V1 0 2 3V

R2 0 2 6.8k



Rd 4 2 .6k

Rs 0 3 1.5k

M1 4 2 3 3 ptype l=1u w=1u 
.model ptype pmos level=2 vto=-1 kp=.111806









.op

.end
