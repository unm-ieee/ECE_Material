XlxV64EB    15d7     890G�"��߽����GS}�o;ȅ�C�v	4��b���:K����l�8�hZ��X�`� �{�U��X�{�G�O���<ra0qK'������v�Z�9��-_Q���/�:w�����ı�BX�M�,]F%_�_y�m[�NF��%����-S�:�w?D�]jч���/ \�� ��²�L��еf	2��U�U��t����S՟��a���O�kș�k��ϴ���E�c��ȜѦ]�m [�xUo��
��g[ª������>%�� Q�}��P�#�+FAl����K��u��!�6�t�p=�Q��E��
�}�L�?�׃J��I�쨿m�����@�!�ܰy5 � ��tse��Y`�l�I)*<��g����x�ww�Ȧ:G���ǔy�� >Nf�{���t�ƕ�����g0�c&�i86���)GqE}+B\�X.�Yn�~���J��F��z}2���x�n�rxvsH�{�<h���¾2br����&�wC\�F��L����Ɣj�&��H=f��j��b��;O�Rr��ﻖe�qV4Y�h�#2��ki]㉕wÉ��C�ܙ	�EJ�1�8��j��K?Wq��m��Z�R�4�Ο���S8>Z��#Q��B.i8p�	���T58={c��'cr�3�� ��n�|_�;�Sf������}����ɲ&2���Yg��K�E�_"����o������8�(� mtP5
��}Y�XʎW�?Y�d]�8��C��h����+��&�6�\X ��j�x�����)1|���(��t��N\��1�y�t��$�VM�Q�z�6/��Y�7�6��ן�@i�p|�/J��W�i�����uJ�
��k�{��rݠ�BqWcW@�a,u[-�T�����C_%�7�YI�����3��P��U?���\��m���j����*y��W����YS�N�$�\XmQE�EG��Tn֎�g��\�F����*��7a	+���Շs瑟��5�����_�Y��W��Sc��;���E����{���#l���O���oA�!t��Z�&�1�֌��r�f����{rZ�?��8d�V�>g%p�J��o�?kˢ&�t�I:��dA
��-��N�XB�X��q��H��	�U��;o\���_F[��\}���~I@�㺅֭���@������eM(4���b���`�W�������
�-���|��W��o�3��V�nm4<ԫ�V��"��<o�w������WY*/ZԌ��ǧx�$��ƭf\�^z{��1.M�
�#�Z0KA��y��� L����!BBK�Q���������H([�t�u�
������G�>�J�b7��2�v�G��7@&(gB�TSD�V�s72E6^�e�U��|�����RV���85�o(�&D <���E�J�O��ɤ]���>�������.6$@�aИ?�Y}?#�ی9����ҝ3�'C�WV|�$̽�Uϖ,���&���* u�����lG�3�����k�b5��H�V�Ğho�W��Ӹ1�
N��c�y�{Ǩ�y% �/�0Òd�
dN�g�������U��w"|�,3���w���f���aI0��[\(�%����cXr6�|K���ɀ�[��BT�y���"oȸDHKY=け�9Ŏf
؟*���_�m���:P��ЈgpQM"$c� B��v�����fV�KΫ+�a��[;R��q��g���J���⒳�
	��	��g���P�������O=
{Yp�	wh�wu#���Z��P��<���[�Ze�`�����4��~`]����q>��빃��o�Y�!�[p����6�Z��8��ؕ7ɟ
��
�LʵkO����ߑ���^����5|����8~��P��.�e�"�����P(5�W��� ~��I��\OR��\��A0àC�$��f�Ș��=!Fy�$0``	3�)y5��v��%mM���#x�9�� {�Ζ����X�.�d��.ت�� ��<;��ȑS��=F�y�.��>����:�~��$_F��8�-�}�3�rMb�o~1# �,/=o��/1�^�f��]�e���{O���"`x���dR=���Uol��\��+2�'��޹~灯nhIs\�o��(.�