XlxV64EB    14bb     820��/Ȍ�҂������&y�����>k^ݐC�?\%��Ǎ�i�ۼSz�}i/ߛ�h�dn�u���P�Ku
�t�j�I6MT~�y��C�}��v( ;���Wi��1d���O��2�h���^�5w�f=;17koǆ	��N�I�}�+�.Ł���^i�DI%�R��~��U�m�be��R��/d�frb��<t�����rN��~S��c�p�W#��֭~ώu�b"�Ճ���zpJ�VR_�"�d�7�S7�E
�������Yvݺ!:V�d[��X}*�*z�Tkr��L;k>�n�� 
8)�Y��|s���N����C<�-�fq���I�M���a~e&v�Q˧Bno�IӔ%OZ���4p;8N��<�▓Y��Ftn�W�" *[��7�Q�*6�g��X����E&�X(����8^��4s/�����И"����0�ˢ,���v�؎�[��=����Ng_
��u�Ғ���:�_���]���?a^W�J�D�c�j��h�'�k�ĩ*��)T��ZߒRV0]�����P�N� -����I+$����P!��Ǎ�l�U\����ǽW�)��Od�@��C��^����0<��!s	�⠎q���C�O{u,��;�-	���^��&\,q���	����,9�
�����I�<�Jh�cQ�?�'�+���m�33P���� ,,2m���p|��ت�3"CW���Zr��7AH>�[����ѣ"i��!2��4{��h}��j45�y<F�&�}�e�RE��K��t��֘�V'�s-e���ۧ�gLN�JS4�w�i�X�d��	x��ɽ�a��R��R���.Ş�QN�Yz5���%0� ɍ̕�grVE��ۂ��T~�e�b�@gu3��u�xW����t�lsLYi���5cd�wb�+��ȡ,�d���J7˛��G�ҷ�Gz���&����+䞹G�J���n���*n�%g��A���Vt��Y��Cd��������u�86/�d��M/��o�����D��̊*�p�����^Y ��Ս���*,�P�W��f���&��n�i��G���X���p3�p��Ո���K	d8�S�ާJ�!r���`�sXFe��!��p#��88���/f�?��S�.�m��l(�n�e�q�;���jo����R��n%kx�Yy.��^��}����!�I<����Q���f<'/�?��u3�wBr��>�^�ʄw;O���16U�b�\q��+�}DU��]���V��?K��]��_�a+��H�M�B�O~U�R(�a#�(�pkP��|�/��!y�C�"H0�>z�g}�-�-�G���㘁�3l�����d�A�Z��I\��evld��Z�I�M�]?�4�V��>w�)
wa��#V�Z�E=��?r'�g"�0}g�M�E����f��3��wj[u��(�[�Fj�ޜ.�o3� /�c��j�B2���XX}@[�a%&G��6�ܸ����ޓL�L�}kcZmW�UW� m/A�8�<&v�-P��>�e��$-�4õG? �s��[l��%Շ��]���{e2p�G8z1�_:��Eٳb�;��w�*��OA1�������kS�m5R�oQ'�OZ���]��V��,�6r���� ����_�2Bt���bJ,�pB�؇�t>L������ٰ����K_Z������"xw����y�S��L;Y9�uPQ�/��~`�W<��I�&fGHc�̋�X�[Gy+xh3�?.5���
:Y4"v��o*yWU�;z;1��&Gj8?�NP����^;����p�q�Arٖ�����n�f�]�k�����s6	w0�D�h��B��� �4Y�2�3���K���5D���<�^�k/��z��Is�X�y�{��/-joY��u^#���G�_�1��7y90��j�#����{�V��~"h�*д��ƅ�N��]m�P��O�`�������MB���U5v�)����խ�=�'XL�����>��q��a���J�0N@/쇉=�F��^`pD�U�l�