XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w^�a	ۛ���mp"�����K�Q��19`����y��qwr�����LG��JؙDg�3�	�d^b4 �������VbO��K8O(,B�Q!R��f�?�L�6UN�@8/�
K��D ){z�xҺ��D2��U�*E�������D	JE[��� �L��3��in`q	���4��i�l�}@��2Kz1�����}�*8LQ�~�����,��M��-A�lB����(x��/���!��h��{ �6���������@G���\���47`��zp���W�]�;�r��p�����2����m[T��Uk<���q�V����^v�D��j["n5�� �zdxM�ۑ�q������ո��rLJ�I����	�s�L��M��������t�,m��~3�A�jj��K�>/q^���-~�"�p.1"�fk����Ƴ�7��)�x�9^TW�P�=�-�9p��t�ի�I�x5�B�/Z�n��k�f�0%T�?[Y��tK1��XDAX$ⶰMZn!U!�ΐ��& �)�k���"r���3˃y̜Q�.��1���hawٵ��
��F���cZ3;�:BcK���N��7Ԛ:��:�	��/��I�C-ޮI��!�D�B���{�`�6ZU� j�f���������!��=B�(΄�	�V�!���,�6�i�ґ�oM8D�X�O�E�1�Q(8��vo'_����~o"L����U��8�ܮ��>�C�N���b��;]�P)9�e��J���YXlxVHYEB     400     200	ညeXb\&J���I��7`AVh�gW�d�~'77@���)ȡ�F��YM�~�V�ZS�/�>cxo����-Q���e�N���J�^��*?]�z��>7�E&���)�^?VԾ��	Ͼ��>!�9����lE����'�?L%����&�G�]A�g8�4#ӈ�$4�x���J���q0o{,�[��4hs�n������(�Dz%Ur��V�P�;�[�Yt�D�0���s�!
Z�\���o���l��#s�!5�D�N�@(��Z�[+���/"?j�Cmb_��(�mY%�._)�H��E��U͌�iZ���h�wJ�@�J5@�����7���S�=�ku���� �'�@��\|BI��.@DH&v_RxhCɾ���h|Chj�g�MCvU7�lXZI6ւ��L���
g�,2dI
�lSV�2A�Nf~���Zw�����MaV��ȪQ������8�5-�dZ��B�K�3DD{�}��?=㵥|d������<��XlxVHYEB     400     240�Vº���~��i`=��d��\��7#�iE,�ຖ�A
����\Q]�I���`��K��J�����WL���e�Lړ���em��n?��D��$ޠ���	,����{DOHʦ���P4c��H��-����yCH_�#��`T�x�_q��Ŷ��&�ܛ�6�Q�����
)~�m�t:%V�����}�pK`\� l)0L���+�zn�ʞ��C\�<��k��i��bt� b�k��ȡS�J�P�l����dN4jp��}��d�*5�Ԋ��E���A�������a�_|٪�:����%�����{�6@gѬ�mL��j�H��)-%Yv��f��x��YD#W�d���B��i�mi�:]_'v��a��5�M=��QwW�Ȇ��I>�6N.���O^%Fh*�Z�RnQ,�S&���39�F׭(��'��m��QU)�H�Hl�`�?��h�e~.�+&��4s�t�M�n$(f��C7+Q(��9�Q�����uu��E���~�����L��߹fq�S����<���?���T�斪���`�h�C}%��pS��8Y%�=Q���4�n�!XlxVHYEB     400     200��V�ե�
�2�&\fh��[�=% T�Q�纪�+�\4��OA�O1���Q3FL����!k<s�Z�Yk�|G�k�/:٬z O� _X�С�hUU!_9�z4IhiQ��H Ó�$&k^���r_�v�Coz� �W�R%��Y���SL�8�ڸz�8V"��'�'@08���/0���*��ũ7qK��g>��]��|�R�d����ψ�r��j�hJrG�D�~�|���r�c�R��`}X���Il�B���q�Ui	O�/Fhz�I����v�S��Á�פ)�"궏��@k+�5�ch�����X:���o��u��i]��Qa�v�����`�e�\�,N���:@+���z�N�S&�����:�a��\�l�o�mY�I���K@g?��eהص�f���f���_�$��d��r��y,L�d���Z��H[����U�o�T�^��``�3�'���2�y�b��&I�5z�$$���V�	後��%���6�2��j�O�RXlxVHYEB     400     180E,�c�V���2��Lt��tL)�u7A�3iu��+��)�甤��ua�9IZ_i�H_)�1a5{�ɍ�]A1W$�A�%Yk���C���	�l��ޑ�qw�J�4��KnJ�X �{��]��12�r����7�oņ`5s0_Œ)~�=����
���<Q����Mm�XwA��s����ڞS ��S>�S�a
$��pV��4U�p�������[� �|�#��Ɲ@5�B#`N\a��=B$*W6"A�ht�#:$�����Bo�;�0C���k3�,������aD,P�LR/�o������H����"�(6��� A��k@*6� =eN3Y�O��֙�ؼ?4{e����#�KQ��pʌ����XlxVHYEB     400     1a0^H
�5OZd��k��G��%�<�YL�����:2�����/�#�\�O����nWGE¹{���so41�0�>�&�u��t���jj���%�]�Ȇp.�0�O���>,[�w��ε���(��\sR^�@B�����`,���R�K�d�Q4��_��N�?q�h.�=BѾ.*w,B�F"gr^0�5x8��%k�B����?;L\�ɢ����h��DM# �♯d
>�Ğ��*�h�{j�����&� P6L�e�K� [I�����#�ʐ�r�0�� U8M�/2���)|u�J�+�"S��6���Ͽ��v�?|�z���Y�?pB�����.$qL��&�����p��Y&�m����aPٍL�?d���gf��{�L���;���u>Y(��>�F��U��3ߢb�Q�*(j6��XlxVHYEB     400     170������Bg�^{�#?�L#�[�_β�BږyL��(׍J����K��	�H^*F�`r�`�	1�Y�Y&���LeRQ��CΝ۳8����*����7"ӱ�t����ʎ)b��XMI�<��f�N���6kY�B�>ScJ�8����t�|��R>��'/D�3�V$]�>z�ם��e�~(��;��2����h�*r��cJyM�ځ�!B����u�4�53psUڛ���qL�7���:�:����%B^�+M"��V�tM$��߳�5����nb�zH��n�i�,�-�,�h9��ݩ���NX����Wƾ�	�b|&��v@��-���o����_�'��l9ލ�����R�9�XlxVHYEB     400     130I�X���+���]��jY�����`���'��vY�].�I|׋�I��ضO�F�"�!#��$T�!1-SX!x�,��f"-t����%1���$�L��]s����3�����ʯ�u����p�v�t7�����8Ì�R:ZJ�>�h��~\�E���;ڒQ�����L�AV��1eq��
�y�o���$Mλ@q�WrX3���A�d(~��o���c�/'m
�?Sx㼙e�G"S�s.D!�aCH��;�$RqR�6�nxA���0!+�U�˖�2ۡ��;�@��7{2��E��XlxVHYEB     400     120@��hF�엯z����mƮ���4��nl2@��w_͖&lc�b[�W{�����z����0@��`��;��A	��B�*f��	~M�\,_�`�q���M����N�W)�?ot�eя:`��n$RU1�@p�l����Ae�P�]�f;cr���FU��tiG@�FT�ǃ��j=�i��&qBd� )*a�y((�P���4�L���ؕ�9^u�����0��1����9�*Ӱ$�k|��o��ĀYȫ��K�!6y�W	�j�d��/z_�9�:O1���j0%��W�7XlxVHYEB     400     130���3,��v=�7�^J��VK�ڼ�u&����ŔЛJ	M�}�Vd��T�н��3c]v��Y�����m�.���J�6�!ts� ��{��
����^�7��9~��vŎ�-�z���eJ�����%9�Z��9v<��G�Ƿ����#g�Bry�Mf��ʮý�d��T��.4�Q��_��r�*G�[^��=�wŷ@�֚6��1��|~��� �ڧX�4�$�9��xm¼��`5'l���sp��0�<V	hզTc�
35@��NM�d]
%�ybO�n9:\O۴����z���8�Knŗ�]8XlxVHYEB     400     130 �?�.�֏	���b�|����c�
�k�`�٧xuo��VH��rP��kJ���>���\����D����ǝ@�U�:r��^��K+Lm�!,�`!���%��� �:��-�9H]�oK熝ƃ�ڼ�6< �e����ݒ�z�]�$b�*��7���q�{:�a����l��}���|\�o���f7B�O	Y_l�;j� �*�Ù����j��;ā�5#|���G�x�#Z]�{4���aӊi�{���:};�e�w�;�-�͔�#^?����X�pX��pL�o�Z�$��y�XlxVHYEB     400     130>+�\�dc*�
)M6f1��F6,�R��i��;��[PR����Fv��;,mC�Ûp��a�:�f��	�����f��
�e���ǀU郻���@Z��ꮅ��m^�56��=k|���>�/�Ϩ�%� q#�v�ث��g�W�L�+s�k J�����':\����ģ�o��J�EMh��~  ͕(`$���O�l��b�a�����|�I��(���z^�}F���34��$0B�:O *�Ɩ!�Ь�E`���f2|&r%3(T��n� ������Фd2��\ʳx:2g*Z�E���6�Ì�"�XlxVHYEB     400     120��C�z4��~��>'U&��a����r�w���uh�n�{@5���T����]&��n<��?�;X�4��\��"��-!)C84��\ $����Y�2$����q�G�;T��t�zu��d�A#�B:��h��\O��Kg�g��$ֺ��}*�a+��I��V�J��x�"�.�!���jd3�Ԍ��b&�k[W�]Ѽ��i�Bʖe9M������G�֋�b�R3�<�u'�Ά�QY������Gf�T{)8����I4K��0.��k�{K�W��
�!O7)0�@�o�XlxVHYEB     400     160X�7?��`�%?X�w\���Q	�r�B�~�}��5?�fY?�Ώh,�c�����P6��p�g�{�Muڜ
z������Q���Ǵ���MԦ��\lW��Q��x�:8uQ���ITA��4������1�s��	��C��M��P|�ó�o-n.�FF�?RW��˞����fU�_�@�y���_�e4z�1/ ��o���r�
?Ʊrl!])M�c�;���H0�P'C��0��k�b Q� ��\�F9b7y�#{̃����;ȋ�Z545���4�F$�g�/��Y�y��RĢ���V(ζ�.��9_rS�	�_�lpdF$l��L�pH���XlxVHYEB     400     1203c������:�v��~�vӪ�H�o�����R^�]��$�c��K���Z��7R-�z+@�B�x[͵a�~�8߻&�{�\]T꣠�rNSem��o#p�n��<�'P����[V�*I�d]��������5Isx��6�(7!��OyR�ƅ�#�[1�v��@]��S&��)�l||A+41 �ᬄ�|g�� a�Bc�x��8:մԲ̶9�R}�tq/��l1�S+�l���#�.�\��'2-׭�����to��^6"1�K�'#�y8�FƜ������eٯ�:XlxVHYEB     400      e0����,[u�Qle���
R{��x���I�is~�X��zD�hL]��=\�������&u��SB��pg���d�a�S����K[t�R���T<۩�Y��{M�C/]��r�"�6�A�;����Nȁxb�����t��ԫk,UP�Q��7׌~e�p/��%i1ezz�P~H��xՕ����d9=��'Qp1���}j��tCOL��<�x����VXlxVHYEB     400      f0��y��Tp/OQ���a�rj��.��{�.���{����v5YQ�Z.�oj�4en���'�Dr��Iu��V��<����[m��?/ι���d3��|�}�g9�x��o�pn{l-oB&S��Ie��>�'�p����2�>o,�١ח�\���p���y~"�|�r_���n�� H�)fѕ��:�F���>�G<QĊ,|�˞�¬�>��돂�e���4�����>i��E~�)�i��XlxVHYEB     400     160�@�0cx��/���@�⬣|�S�1hZ_7Hǜq\�?�V/U�Lb��3��)�+���Ӏ���!\L�	�h�xFX���)�8_�	�B_9�'\U�vҲL��e�Ř��xۢ��,�{Uf�;��JV1�#�l�H�Af�SBH�9|�1lS����;¯[�=dÆz�ۄ(�@7�@��ٞ���=±-��h�� !z`��24���Ӊ�E8f�|�VÃ=¢Ї�-+�����@_>Iu*�5�Qc�L57	��+7��m,y��Q���
Qn�˃�.ߢw?�m��_���v�R�}0[�	�tJ��T���9#�c����dXlxVHYEB     400     140,�zA�'D���aU���7�������T��>�6�N�%��	s������P�)_#p9���x?Y�k��jC�E�j�p�g�Q���ՏN"0)Ƿ�$�q5
`Z��W�{`�oЊ�A��z��Ő9�B�Q,V ��rH���m-�����L�E�����A�Ny�WYɈH�Q����C	�8��AZ;F�O�j ;d�V@�č`.�lpa�׋1�v"0��!���Mҩ�`�� G���5EB��T8�6���U�gӣ�MzH��A��Z���;�������g�S.�0�&[赜�.�x�����B0���0SJXlxVHYEB     400     130��٦��Ew���/&:T��i����;�>���W\�$[�߯�'�0'�q�{�D��������.����e-�2諦�E�f{�al�e9di������LO��J��������Y~9w�#*+����ܣy�%:I|
�sڝ<%o���I�>������
��D����5��ES����Ot䞰I�(�Q� ?^�u$���|gC>Y�i����$HI�5�i,���~"���p錟ny!�NaR���>�ߠe�;e6�&����"�V_bGNy7t��P�x>�؂�HM&����l���XlxVHYEB     400     160�-��*Y��P��X̪��:
�^���ɵv�06[8����XBk��P��'�v����%�.��}��	;�C!ȹ�G���K��13���,`�a�t���*���0'�������
�4T�-�j
m�M[x���o��m:v��~�Q")��)�Q�{y����J~W9F���R�'������r䨇�Ͷ��)�m�~�	��M��A( �w���/���MSx�	��D�Ơr�c!R�&�2/�&<���)�]�i�Ɩԝ/���&[�"�Q^&gu�|*)��]&=������aM�DtI�@�˗�ޙ]��� ȿ1�K�P��_i��ـ ��r;�{`kZXlxVHYEB     400     170,��^�n�s�h/ql N�JђVA�\�x���:�_�]���T|YM�z���*��:qѧV�4}���xFZ�3~���C��>ޜ
c��8yEP(ia����%d�6-�$��G�BX�Ϯ,�
����
0�$�D 䢪������>Ϗ��&k6�j.��)[NE�i,�ȏr���x��)0~�Z�J�
W��#�T{{�B< �Iz�V���hdf�b�l���Yќ��27���E�d��l氥��s�ί��{�5I�G���f�c ����u�VǮ��Y|+��g�tOMt�Zn�����إ�J���Aݏ=gC�);���1��/��9��֔8�[N�(�q�v	k��f-������TXlxVHYEB     400      f0TH=�y��\l�/?��ă%9��	��� � ��qo-�T��v�T3�R�!�aG�u�Rw�P=K�FFDL�ꇦv�����N�gt��v�@���/����c��!�с��4�w�X^��(���'��qb���OT�	G��.�墺�I�4�����ڈv v�yfz����4]d��y�F�е�w��\yu�FK9���j�򀜈��~+�u2���?�M�sd��K���))tq�XlxVHYEB     400     110��q��AH���j���Qh[Я8V}S��E�]� �B����Xٗ����&lc��]�āWؒ���Q�"��lr�J��W�"���N`�S��y�b�ˑ�h����7��V�7bIR�oO�����G�
S����a�F{RDW��M����˛��n� f
�ͼ��	�c�o��,����a�	�
�t�:��sW4�溼j%��+�e���*�[����܋�w`i���:@k�����B���bT4}� ��LA�.XlxVHYEB     400     140Z�\�ה�g��v{|�_����}��� c�b�a��ue������Vo�Ma��{"�\�z����k˭��
�FI�A�N�?3Oes���+�-cA��cZ��ʉYq��w�OQ�;�[`����>���Os���IJ����!�F(r�F7��u�h��8db5�~W,:�ͤ�����o5%Y}��zQ~M��^��u�o%;���u��b�(�n>'@IH?��3����?&�hB��~TN���e�됃"�F�	�P�!���q�M��S�{'�Yy�j>x�����X���l^i��A/C�m�/XlxVHYEB     400     140\��!�`-�K(�4�w��ܰޕW�ru)]*~p�0Ҙ$���G9��=1�y&o�~������l���oWb����`�i�˖� �+�2����/�J|Fx��[��-
�<�j�	��>����]�QE�%����I��@Z���Mj���4�� Z#�שi6�0�eCl�GO�+�R���3s�3z���a���w�8R[�v7&�Σ���-�1��[s��F�q��p���.���"��< �()AD�1�z#\M�;��<��|�3Z�W\�{�Hw+����}�� Y��Đ5�$�) � w��'�`�QXlxVHYEB     400     120B	���3(ؔ�-,i3.`2ȡ�zt��<�x�0bVh�(�QT��+%=�Z��q�%L�`�%����YK���N����ZÌˋ�T��Rt �3����DOD������c�>������)�o��!�Q�G�j,@����TA�ۄFa��|���y|��y�I�����#ٴ{�n�/�o;W��0�>��"8X6IG��f�Ԙ������I�+�J<�kN�񯐵����"�.�ex��/L�:D�&�����Ӹ:9��t��qʘ2��{�WpO�ȷ��+�����)XlxVHYEB     400      f0�
��x+��nS�
?�����9���ɤD)IS�7��J���O-=T]��6�I�=#�e�̄�������MQD/�F�8er���3��Z�ҷ��+Hη�����ھ�Zj$P�R�$#��F�m4��%k�:(ƥ(��^C�߈ob&�"���;cT:=�����T(gX��!E{�4lt�����8���Y_���}���>C�1�R�H�d���t��;���Iwt�`p�*XlxVHYEB     400     1303�&���y?V���oT\aD38a�=ڼ�NVl�8jds컌�#g�c���\3ڄ^����\�`�y~�ٖe>�Vh�GO��0l��0��R� �!/�;E��|���k�!�2��`�M�/g�� �3T�yC˛.:�����[�7��JI��PE��E��u+鿣3���l����������z1�֙�E����O�}�[�H�>--q1��2�l�g����a"Z�k�HSN�bf�،�io/��~T����E��lj��:q�+[j�9nۚ2�)��6�RM�fvV��x�1t|XlxVHYEB     400      c0��7�ìo����oغX2l�5���L)���U�A�� �x[p�d)�)��՘�n'=T6��,��ƥ�N(р����8�O�8�^�8l��u-�+E }_�Ŷ�"�oV���v�-���phc�-'f����A���v����]T�,�Nx%5�z5�aJ7�$���t�mu`Z�d%$�X^�'��Qr�H�����!XlxVHYEB     400      c0Eq��3�C|-�Y�ף�&��
�Y��	�g�[� �6����
 9��]�F��ڋ �����ן�����"	5]��p�]���$*p���u�h�����D���K��0��`��+H�7�Hi��&�4�1�}���Ǉ�N�Z�؛'(\�y�a� �������4��:�{.�B e��m��K%�̈XlxVHYEB     400     140��l�]`P!f���#�u�oo
�n���)R��8��O�ڽD��Z��-������O��$��V�UxԌU+R(
��� R�Sf�\A��,S�+��7����'Mـv�2�(�l�
_�;v%I�|e</��`���Nu�Y� ��y�\���2��)n17��\s�8��������Ռ���q���t�icޡ�S�
�����C*�v���h��!R���=�aA3�5�;/�P�o�kf�s����QBA��1�U��2MKobm��!��Z�����O�薆.��;ej�k��|�#r��^�y$H��=���)X�1�2�XlxVHYEB     400     100�YN T��5�F Q�B�C��7i��N;�o�FqU#ٰ�08����l����|�&c�������t~�%�%��	��]��c?R�V�Ƙ;Ol^uj�,e�b9��|����5��}5�$�F�v�Y��{����m����;`|�Sng��󮂢mSF���bI��	�n}�d#�	��ptG�q���^�F��&WU�a���$�~�D@C�U�c�zOMQ9�(*�+�<u\�R�l��⢙�J,�@�
.��XlxVHYEB     400     140Xf.�.�a�d�{�B*Fd���5U`�&�9���&�8��%�9wL�rJd%�����7tztNyy�޶1���)����{f�T5J�`a�NNƌ9��,�4�$�xf�J4���=�����e#�|JU%g~Or�V�.^zf!q����<�;A�>Ţ̄ݳ��?��-�`���Ƴ��|����d
�� �ڥ��sڄsdR� ��� �������.�T
U�mG&�+^�{-ȳ�L��7���[��/�BK��/�9���K���1����$��QyN)����z���6�!(�ePۃ���8�M��b��,��M�v�P�fb'AXlxVHYEB     400     140 ي��!:1��}�����Iv���N���J$������2q���Dww�ׯ.�f�(
��0��n�e�C%����[�!9XT���xH��Z���g���������e�	���l���B��Br�\8h)0�cE���R9_�����(���2���9M��j}_<�'��		mp���
�be]��C*$��B�o- �# ��qT�&j��`i����`zYiS����u�o�S�_\h��娭��8(���k�Μ?di�0�w���<U8���4Lm&�Di���R�$�[˴ӕ;�G׆��f܄A�A؝0j�~����XlxVHYEB     400     130h)2p-�)���H�j2x�Cvݽ!�d6��<LW̘M��ڛ�<_�k3�E���o>�����7���N��a��EEL�����*���M�$���I�ID��dY���3�nx�1�
��)x>뵸[&�"E129���޴(�A�!AZ�qRfhDg>���%��I��~MS��v����xt��-��P�U��a�UN>��Mʥ�	]c��nV�������"%��9F[����%T�����M��Ѱ���Ll�V������"Dֳ\�c�sU�{N.���b��'Kpu�ʣP�xqN��C���#�XlxVHYEB     400     100#ṷD��a陠t�y�Z1�`���n���b'�a��c�DY����M�Fiq@Ř��H�xm`Z]H_D2i���������y X���z{�9ک�G�C[�6lY�yͷqH���g��`\�-qpH�&�BR��{-Q�l�)V9l0����|A�/�4X��V{<�F�J��Qܦ�.,����)RS��[dZWc.��j�ON<�G��cZ{U����07�s�a3+qo}{�HZ[@�v�r C��8��B�tXlxVHYEB     400     110qx�Rg�gkjǽ��_9܀�}��>��/_q�(�v�2�KG�[�Y����_�{w �&W�U���@fyz2w��^�63YY�8%��x�	Y��mR)NX�2�(|\$�ۍ.�1fb�[�P�3�-l	����x|��==
��}��p_'h�i��T���P�@��yԡ6�l�|���h)��Ȅ�.]:��`2g�_::WT]0P��̟��x���$�*�\�-#oB4m���f�w���b��"K̍v��f���#��A��j�v�w�ҭ�IkXlxVHYEB     400     100�vb	����l$e5D����ix#���y
'ou���T�	}����\�g������n&�Ѧ;,�p��\M&�m��%�T�0��B~�o�3I=�&��P�2�*�@����c�`��r��ʌ�(�D=�4Y�|��m𖷡�+��!���� ��|�}qR���Ū �-޲;r�[o�C��JN��l+�*��KN�+k�\v�=�9�����M��jԌE'h�'�P�(��Yr@4m~��ݎa��������KXlxVHYEB     400     110ɻ��
��׻h�� /�e�����ݴ������p���)n�/\Ht�&c��-Fq��
w�;_�Nx WM[�_������2�gԼ�>�T2�B�k�X���o�"'{[��DW�	*d�d��������_�?���Ƞ�(�r����(}�K87[����AG6�[{�Q|q���@���ao�����G}���#K��P��n��c�tnw �)��:[��G�=	��8
)�=��%���e��#�W���Fڥ�뚪��n2XlxVHYEB     400     110,J�S0WG��=@�O��	�&��a|�i��M,w�+xfFq^7S���Č��9�4�ځ�t��;��=���Ud�~V"ӆ/1p uuM�%�g�n�{���؎.���a5�d�(�#U���r6	�T"V~S��^��E�K�P���SfӶr2��
g� RX�V|�l��C�|HzS	r��]3u�N���i3Lױ�3�@�gi���'H�Wj�q3Q4Jߴ�y��}>�f��[g�\2`�@1Fe�[���h`H0��^FXlxVHYEB     400     150��3K��>��XD$O�l ��n�{n��ߤ(��&�}��<�N�w��0o�n#J{]�=|�~�Gօ�����t���H��鰣)�UA);ƋRǝ�ȣ=Ho�L�.��Vy�De�彜Sa�����d�C��D�!⟣ޯ�p�6�(FZOH���F�3_Ky�Wji�zo��Y��Z��Bj�c?f?RCɄ�s�+3���N��-���$�n��� �~jE6*�^�q��[�]�Ͱ�5w{��:jF��(Ϸs8���h�����rg����J�����Ԧz�C
��8��<��͜Wm��XN�*�փ0��"$ɉ8�RΜXlxVHYEB     400     130��� L�h]|�� l'"���i�8��p �+HS6�-xG	
���~E��Gw��4��5��F��lr`1	QUyEJ@Xֶ�'���㛩�>��5�@�ע�9Ma2��.��uM��r��ps�5ہ�^��k��2�8İ��-�~o����}p�;cܩ�-�$��2��}0��0�7}��	�c�D�᳝K�֯�W��9E��+���2�N����������_	���E�D��3��.מ�`��ydrx� �ݚ���`�]�9a�0���,S�bNVh�Q��� ��W�F	�XlxVHYEB     400     110ݠ0SJʿ�Q2(�Sqg=��`�=O�
v�����tzq��v�&�>\_n	��-)a�(�>�yoPDQ�l��Vg�0ꛈ7]��+�g�ɟJ���e�0Ц�&�'���Bh��R���q�0I c.���]�x}�������=�Y�V�u��;�S@z�������j~t�\jQ��W�&DZ���������.jK�*��M�#�
�"-C�gN�w:�6��Ք�y��v̭� �g"iu�7��j���a^6�Fˡ�#���d�<[�M�QEΎ�W�XlxVHYEB     400     1b0�w�e�c���r��>(��xR�q��1���ª]�q��5+�"_�<�vB��78����x(��!$I�Uf+[X� �Q�%��6c����|bU�U^~2�����>6���Q�7����a5f}@�S��'�cg�(R�}i�Ѕ/����������d�jJ��a�K.)����'�f����:�C�ˤq��y��˨�,;��K|���e��(9����O�����HI�W!�?fz���z�)���N��EI����a�ܜc�h�� �����1���.�	�{������Cu�̨�!ǫR�m>F����O1�܄����O� $l�h�9��O�h�b~D�W.����K͡��Xh��H�+�:�m��^E��O�R�X�
��d�� ν��ݹ�Y��v]���?���p���Y�w��a�?����p0�FXlxVHYEB     400     1a0�y�	�$��1��L����&7��*�9X����R�c�7ÿ���n�|B�3�{�g��?l>�?��}[��K�(ތ:��G�˒n>�z���l���ځ�Y��-���g��Ӌ�1%�o�YW��e���偙�5n��9��!�;�p�b�a=�A_��2������e#a������i�K�5�l���s��wf޼�s�TV:�Ӝ�'(��p(����V���%���!Ox���;auN��b��\��&�uF��g�Y2C�bT����Rm�d)����vf|x�Qؔ�o�L�GÓ�6����x@H"Ei��f<�H��"�_A#��������s�0����'h�E-s�\�=d��UFK�i�=C���/;�I����6�Ɓ��\v�v��B��]C��[��:�XlxVHYEB     400     140讨����v��5��^5��澆��o:��>d�AT��=vؗ�A�i��w�C�������A���j�I]г]�`(�y��B�@Հw��g�e5Hg�¨�s�XȠ:p*j��� ����m�����aW�A��P����ġD¤����X���Trպ�D����?�����1'�� n��)�ýN�(*բӠ��<�~����\�b��h�@WD�9ʕ$q�?�v�~�Tn��z�Ri0�B�
�2X9���P�h�8��cA�f�s"֚5�퇟�ӌ���e��9�
s	�!�|���x_*4��tWwZ	XlxVHYEB     400     150�P���Z��DoR��G�C#[J6�p_tf�c�R㣭��X�p��/ᓶ�۟�b�n�A�̉�{l�����/F��y�VZ�D�q����/tyʚPF�B����J��l������$$t7s��,�p5���q2�:�h?<]�]�~s��-K<u��n�v�&��%�.���R���>,4;C��F}�hu�_�A(��
p��������^H~�)�a�*ʐ��� L��뎵֠�;�h��7��y4p����\�~ͨ�Fvͺ�V�L(�7>FU3���{��V�Ŝu������v
`<?�=�C%B�nH�E���bㄛ����Լ�67XlxVHYEB     400     190PA��O�$�cv�w��q���D��0g�$xA0z��tǐB��G�:�w�y\t_�o[W.q[��R�����!��X"O��6�:6�#��(^}?������݂��!���Ν{m~C5=>\M�
>���{�%:w��/�� 2�H'_�L- |u�Nb�)�ו���x�{��O�Y�K<B�2��P����7@��&���2`�j9��Ce�� ��� �����s+?��4��,�Ax�B� Qx�����SЩ��[Q9��c��L7=g��΋\��&����R;�t��D s�R��@�_L�z���G�+vk��t��.���Nzc�!�u��"�^l���@I�T��Ǘ���a��=��~`�`Tq�0���`>/=K�p�&.>~�'� {���܊�TD XlxVHYEB     400     1b0{���c��i
�jOͽ�̿�B���So�b�A� ȸL{ﮐ��g���� �~?�/��N���\	�ň���SV�Pi�O��� qj��jl�GK�yL�w�Z�������S�.�uJUF�C�nӴ�r��gQ�^IsT��3��r�2L�G� c�� -0�0��82,}��eYy��Av��� WZ~$p�9
�btx�6C�?�]~��?���ǻ�<����s���u�A|��S�PС�^�E��WC�]���v���̮�*�ŃD�2���x����}Pa�Mo�Z���Y�4U3�Z$2[��w/��4���t'�ʼ�4T�����2�{X�6��r#�=C6�c���3:
�d����F	�~���slϼظ��5����k�@´�:���Sh�+��@1�lL�k����ם�K���p���A)XlxVHYEB     400     180�s���x��nf��{~,T1���h��N)P�s�� �A�GOß�zDEw{�A�,��g��:m�,v0U���Z=O΢%���*�&(�G.�SF�mS����O���c��@�g$�N����E�Y��o���8����Т2���ޯ��)7��4ޫ�m��]��ߠ~�n��ݝ{�[=�VZ�Q�$oL�<�$�����L�*mx��2}�Jk9�hvY���얲��<=E��;j��~�p�.��{�Rsa�F>˪����+��>�ui
�2�#Y,\��K�ᬙԗ�t/��u��̹y�ʴ?�~l����;����#n�S���t+�#�����-H�����F���MD|��{�̥��*m�)��M�� 练�������T��q�XlxVHYEB     400     120��j��9���]�v��;�����O��=a��}��D��L�8A-������l���,�@��/�
$��U1�ҁ;��	����:J���]�0�z�?�K8f>ZTr*~����\�ǫ%�*a�\��s����m���.x�̲-�J�0��э�B���ӥ���]���E-�ϖ��y0[��o�	�.C�0�.r���a�#r��RlI�q�d�}@�+%�δ��8(�:��(�ms�a�n�GT��0o0_��*?�}�a���$HXu=n�a�d�2L��z'L��XlxVHYEB     400      c0TsUB�/%�Fj�$KE��"�b�⺻˛a=��#��A�)�����~B���؜x����s"S[,�ٛ�B_y�bQ���M�z�ZF�L�2{�eS�
a�G����w$6��	�i���S)P�M�칂�7�6�ߩ��}�Ձ��)G���g"�)��u��C[�~�)0n}ܥڰ��q�TDG*&6��#�VXlxVHYEB     400     190�藩[2S8�"_T���^Et_���q2��V�K�!1ԷB��H����ZPk���i���t
P��	:�V�o2����&>��kP��i<��,���W�p!���ƺ�Q��{IҤ��
�*�yC!�w�������([��Q*�P?�e����Z�aB�s�@xp�=@�^��Lh�O$���S'Kaa�kb�_g���~ꏣa��r^�R�'��_ ����+5`�֮!�@>� _7٣M�M�G�?W�����=�
��2��Zh��-��A�<��V�U
�@/���A*g@�HP+�?�+��/GՇa���l������ȴ�'B[ӌe��ԅ��.���^�yAW�Sb��U�
������������l�y�9����ޗ��R�v�K�\XlxVHYEB     283     100;�j.Nn����u�c�ؖy=2��6XGY�u�$ s>��_�`K�m]�����p��J�H08k
�����-q�覗�_�R�2�!���ϖ�+u#%���֫X��6`�������1>�wi��.���1�'��?q�y�2/��T�=Li�~*|��$���r_�	������D����Զ�+�/�f(�ԓ�vx0���s��Ea.���:��Ǧ�թ��%�d=FI3��L$f�"p���)�!a󸳗�	��q