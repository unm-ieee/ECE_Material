XlxV64EB    1bce     970c2�(�����ۄ�sl��L�\�45U�x��+q������y�4QU������c��Jy�s_f&�y��<UJr�K�+�L��(�Y�%%�H�u�ȡXRjN����Պs�� ��O�	jGF	�!�󝣌��v��30�4��J}������	��i	�Y4Z6$��)�<wA�0$l�)ܪ���Zk݅U�#<�2^3�S�?.��(�*�k\~F�_E�U���|�6��M��Z��,�����\l�3&�m(�a��䥺�'����b��6H��~'���O�;�ri�cS�/��
M(ۃ��/�-����Y����'��0�$F���&�������յ��r*����t�6^4%|���r	I83�Z�Js�����ӻr�9b}�c��S�'�PI#�!�nxy�&F��.��4M�<S6�-+B�^!\L����(��fEw� ��X���?����W86�L�(fU{|2j8���O�9��}����r9/��_<�Nj]�r�G�$y��+�=k#��g��P�k���pB�9z�F,��-���6�y�]��S����B���6�U>�q�kE>s��ѳ�0��g\��bЪ��ر)?��\c�-��_tJ������/�q��a3T=R���P�+�D)���0��*��Ϭ��j��B��d����)�F65�G�2�׺#�5�(��՝)��L�ˍ�ǚs[����6�t!XK9�Ս=U)<uF����պ!: ��b����O}���qA��6ڧ��z��!�3P%�<P��k�_F�MN-*2���6ٹK�������N��,���u>br�j:���A!���3p��nrZf3	�
�"�}�~��YЉ��YUtZ��Xz)@�(Y��bs�d?"0�-̘�ۆ?˓�K�#�Nl����J	/�G]�>ݻ���Ŝ��j��
���r*������y�+���8��e��Z�8L�%�n���5L� S-���!Oo��h<<��E�HF��G�C���Ø|U�ɳ���Q�,�L��P���)~ƛs�ϥx(V?Z���6"_{�d��Ս�s�X�FG�����F��(I�	�_O�J��V��%���e�}�O��Y���Bv�w4�B�#�{D��6��z���Z�UH3c���S�O�5[������5���V�yǟ��������'.�r�^�F���va�Ғ�ɣeZ���vm�g��2i����,g˳)Q��>+�)`[N�N;Vl������lܓ�Ƃ�q�(�,+p�w�ɪ�N|�:�e��wǒ�):�i�ih�N�a���򙏘�Z+މ��`��ԥ����ᰳ&P 5ۦ��F}L�X�i�G3,I����sp#v�0�ԋRh 
���+,�m��TSn��PTpt�%�v�;�o�/�HA��9��Kɻ��S��o���o/�p=R*52��A�P?AL��6f*��V�m�?�i��aJyqE�V�r8�Kv�!W�g��+����'�O,��݊Y����{� t=�����eqBg�x�]գC����|�,�r�.���UG#��q|��}�P���4�j������x���Ϥ��ۄv^�8V�$8�����G �}���X�)޺��lZl��MQl�d5j(q�3X`�'6BKaj��`J�J�C�t�R���{��tq4q2�<>�[$�~�*�="����F����Ʉ�~��w���uߔ��I)x���k�m�[Q�l\�=���NV[�!36g�+��
�_ל������)�`���cI���2�{��B�A�8� � ��Zd������Asgy�~c����PQӝ��247�ͬs�t]s5��#�~}i,#W�6�a�tH8��	qFo�khҖU�ŋ�p��
��f��jr�e53�`9|~�'�ؑ���4�&�8f��-�7����©���OC�`j��/$���K ʔ�y��ʌJ'ˢWw|��O�0��U�������vo
�Sה��N��c�U6J���d��}��g�L�l#*O�|-ښ������2�V�qȼ��D�U�߰,�qab�TLڀbx�ѐ� ��2���ܫU�E�9���Y�"�+�,W�
����PmǮ����Ȩ���NX�*��^�nnU���/J�	v9�ٿ�mdko)3Z��m-�6��P��\�0_"��2V�u����Z���~Z�P��+d,�S��^q.VERv�$~�Eh��:O���"���۴ۇ��Gi+E��W��B(��������\�6)3">�y.sŤ��E�+�A�5�T!��*�V}��+wŹk�u�����3��Nj���υ:������	[3�M�<s�J?�6E�ݡ8q�1�-Cw������]��+�ݭ�)7o�ƥ������o ���