XlxV64EB    2764     af0.3h�I^U�< vǱ�{�VF6�M/���@��D��2�k˵�r�Oz+sJw���x+-Pw���0CB�&��U��#>�C ��^@�8L|S�p�3�`���Ȼ���:	~�cә[-�.M��'�	T�J�Ⓥ�Z������y�w�K)�����mP������n�i<n�qǆf��w;�4�1'V��M�3aa��_f[����H�G"a�+}H%�;&����ѽxS"�=lb��	M�7��A�"�vE�������d%[(v������D�����_��lq�4F��)�09�zUޥ�QLlr�C���c;ᠥ�e�{�fI�2S���M���	����M������$b��$�(B�i�Z�aX3�0�v�{K��`�9*�^��I��Ȁw�����&:G�LI�0�/��r;(��a.C�^��g�TQE�FJ@���H�ӵ�{��ֺ���o6��1bT�<��(�c�|�yx�����+!� 1K�Jm����V���5��,f�ی�]��Mۅ�QeԎ�88��u�b�x����z��۱�_�"#�f�湣Q'�ѐIt0�	�AE[�	oMʓㄒ�M ���ֿm��_3�7�B�N9X��!�4ڰY��_ў5���&�� ��K���H��.>Q� ��Lc�
rW���4�.����azK3��r�'�kg�rٹ�/%Y��	�\�@͜��>/,���[3Um���U�?�x�0�����ܲ��`л�LQX=��Z�笽@Ao���˥y����7;J&���䞼m����i����}������J�;Eǝ���.�tMfm����G��c>�O�f��B���n�K��}܁Х�F����h����];[ �p�v�'� ��bj���a6g\�H��Ec̕x������K6�'������f���8`�	��L��½+z�
#$�윪10(4Rt,��	.�4��R��q	��䄔M�0-q�v1U���p>�i0Z�oXR����"&iH�	).���,&�Q7vX��oM�� \`��E0�+kI��&A�7�WѾ�Mn?���A���JN^(AD�q��ipJa!���g7w������`�Jk��f�"nZH���w�&\���\���=
^�	kR�C>���N�:�O(	1 �	Uhm�w������2hd>m?9��#^��ƅ��eP�g ?[լ3�������YM\������m�H�� &��xr!�0ZzV���S1b�ݚ[5��2������l>Ipn��:����N�<���:l1;K��"��E�~�q�H�)r��Yɫ��燯8�&s�!���*�Ě[������Pr�#����� ]���:�=����gn������񤲩��UAA�k����w݆�to�PQ�:�^2�/!�KK�֬F���2�\c��yh�|�0]d4�sq}CE�'�����e$B�:'7�
���	V��bkL�ؕz_���#\w�� ������sX���l�gw*>8t'�`Z��w<���J�N�g�@��2;�6}��"?Ga�p��Gn��@N43��)x���}۳ �K��k��")�_������k\,XO4mi�� ��T�j~���<�ƮS��߬s?FXǗ�q-e�a0֤� @����H���u8��v�m4T����u�e��������[���8���C��DP��1fK�w��P��� �s�������g$ô{��k��˴# �}��Q�r�8T"��nsl�m���5�~� sT"����,�U�;e�Ⱥ�W�A�q+��QG���h�%�5U�}�jE	����v�д���@�Q���%����.�D�?��l!�b����Z��t��P������8�up�}���0�dM\�3��?Y�2Hw*A�2���h�h|���#�� }��?#�� ���E�Nx����;�O�z��ٹ*�)!�B�}�-�#j�����ѱQj�(���],q��(�t;����i����VW,�u�|�k5��85�}2�`��p48g��eu���S/��ރaumzB�|ac�%=��� ��3��y�UB+�h8��v9��mVϼhDP�Y��Ġ9$�5��Q�ǪkY�!��z�\�fY�#G/HM�_� ge&R-7�Y�`�"��aUo����{�L���𰁒P(0Bo*,$��cx�|SL�K��~�����W�=�o+�ު�ul��܇�ݙ�	�4�L��4^W�f��{��o�V<ڒ&�H��ls���Ӆ�M���C��j^gh�{���4��La��Ӳ�4�>ؓ'��
�z�u�������J��x��|bꀍ�b��Cw�����??��[�'�H7�h�tl�"��������#�,c���Ͻ��*	��7Q\,�<�U��������@6��g���ċ������s�a�ZaU?��(۫�Gm�ޙy����r����~�ն��'0�]��(]b�G<+s�Ȧ����WKA8z��B))2����}��S�*�8O�k�	:�@�����W��nĨ/�攳���5F�0��d9��x+J���fd`��zF���p_)�W�ͦ���od|��U�_ȏU�����x�"E#%&0��G�ũx�b̧c37����6o��e�EE�=G�\!�]K����w�䤄�I��1�.V�XX�Ҫ*�}ԅ���E�����Wr�;��b���ྙ���K1&��b�h�