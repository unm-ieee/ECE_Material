XlxV64EB    179d     880���'N����UOR��3�=b�^:L��ܻ=�%�Y�U�+�t����Uk5sh�i�?h�'�u��b�aj������c���ʽ4�!A_���O�'�'Rd���3���$��}�c��:��d�{描^+|�� �[x
M���6�d�#��=�B�g�P�nXxZރJɊ:�0����̓���W�p��1��lif Xj��~6G�8�eg]m%@{9�lA8i�& �|�8JG���~{�)z>ų��D���op����O�jF�!��x��ն|;�?H�s���V�a7H�(�K<BȢc �O�j߲s�&�(m\��bc���,Q�� �d�ke�{H���%m���4Ϧ8I��x��5r=
Yd	�r���|-���3�Iq�-ѕt�QJ�Z�/�ӽ 0G"�:�M��tp-�Z.�tr�İ�����]�a_�A�Ts�Lf�>s��eCdX��z�&�V���[VU���~��8QAO��̠��Z���Zh5���]6�kT.�W����߰_v�g)�����\T6�4	<�}�i?	�Rى]i���:^z��\;�+i99��DR��د�9�%���D�߰+u��6^��#P|Q���G(�%���[�ö+�Фt�� ����=Dچ����'Tp�ђM��X�T�U�u�`��l!�_)d�L�5`jL��v��F�����##�3�Ky	N��:���WOe؜K��c�.)�����s�
^@}hG��Y�똺�N�=�L��'ߑ������{�2��:匳�*ǃ�x���_sER��S�`�p�xj�X��`����l�R�|�IA�6=� ƀ>���d�( )��� Gh�gk��8�g��}Hh4a}y��9����a�a�a�s�5���$�\W���Eԧso�ͼ;�ao�d9�Z@�4��A�GA�:���%�Σ�7�Q�����8�Cرk���y{�S�r8���"�?EC%5�%|_��9:�D�b���`��o4'[�
 �NI��M�³���غC�9T f�[(�7�qa�KB�U��-	���~@6[L]-�1�������gM�~vd9�����>f�ULm<90���q�<�N|�(�>*�יm}����sqy��[�?�s�������u¿x;��ƥ��c8{�U���3���dM@��"H���0[�`�Z��7�$-�l�Gh�{z����ඇ�BU��y�[�d��8�{�ߛ�����OY�Y��	�m:R̚:�A�gt�*Wsv�è�d
�f���";��驱[�k7���08���VB���"t}�T�$���J�����Tʂ>5�'eZ�l��5��p%��}ܕ��d�*�� �xRT^�����r-�8'��!fhn@�:Rǧ������z+��'\a�6��ő�n4m���~�O7���W�]m�Kpr��*��õg�� ��5Cg�� D��mŒBS<N\��l�R����PK�3N�F�D�y:S�=cZ�ߣ���5[��6*�Ih�f �xqU%��g5#26)�e�]"�<����ʳ@r�[F�f���.��3OGe'!�޸y)��ы�k����FgP���ԨX��������SJ�Y�	�`kª��ݢ�� +$����E�X�"h,1��*�u���y�l���_	���f����u!����|d)��qmN�Y����_��M�Qs���`{d�6_�g1-�is˩���iv,�d(�ûPdI��&~����k��f���/���[/-X2pq�y�G��a���EV>n�_�J2Ջ�X�N���N�e�����k�N�vl��э� ؑ��^�Z�zOy�hSa��M���\�X�zI�u<������oy�ѩe~�8]*���QY�D����̷��?��uڗ���� 8{45
���;��j�໐�Rf��w�:�Qz��]"O�������� ���Q�ʍ��㞝��v�6��
A�2���N Rn��d�bRO��YÎMm�?[��<��ȍ�V���TZ�%�e]���x��6>Uo��֋�رQӳ� �}���4hgl���AK�����b�-ݸR��~"7��E��O_���q,��eT/�sR.�y]ҵC0�ծ3̃�;*{o���r�wCV