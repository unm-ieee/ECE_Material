XlxV64EB    130b     7c0�t�ᬷ�����%�.t���c���J2�T
�q ���aϭI�5ܪa�Fp����P㥂�6�$�AU�k����eD����9�wuX{",�u(��t�Wy���P��4�r�xO���h"�hIp��-ND�ey�d�E�5ߏڮ?�l���H����B ҇�����ID�U���/�x`x����A�ނ�4���e��\T���e�t0�+U`�u~�)Tӡ/k@+ʹƄ����$i:���ʸ[C �|	d�u>���S@�����.��,�j� (�Z�p-���M���YG7 �$�{�-J��B�lz
wZ����R29��q���t$LMo�.y�İɗ߾�:�fn��2����] t$-�4:��/�]D�Mo��:�|�C�U��6���߂���)�T���͘ƾ��*?��6��$���%cm�� �x���6 �/��-I8,�/u(�����nZ^��7mH1���� Q�GP�(�_�a��Y�(��Kd|I@"�:�x�H,^m���7�̼t�{��E-`���0pI>�Oe+�ѧ\Eu@=l�D��`7�����G�W���(hDW{�Y}�o���AZ�z,�|�Aj )Pod��Ĕ�ّ	ԅZm���	y*(>q�FJ7`u;�-�`P2����Ʋ3�j�d~X;�4�a,����$��*6
�G�K���R�~��Ғ�<�(�����9,�}))II\���vy3�bo����q|j�턎���4�8�ZU�E�p��5��}��Go�|$4q�)&�Xd| �"ͽH*˓�G4�ub�7uz�9��aXK�b�>�!���![GT.��71*d��8mA�B1���S�b}SϷ�n7F�����D��q?��Z~s1A�'���h/�Y �6�+���;�|�8��J���O�"\��n���!V@�3�Z�\=P���	��>�����i@��G��k[�����:<��"��Z�=�k���3��2�˘��A�&�,<��E���|[t�H_ϳ'Qk-鈅*x��+l�D��!]��x4^<f����ȼ��Cx��@u,��N�ō���]�1�N@ r-48@� �T~5�*��E �n�����Bh��M���e�z��۹UEQ0y;��5��@1O�V)��"oSVʍ�ub����A<p��rc����ӻM��vPj���$���ux�t�`�NӶ�2��ma�������I�۰��KDXv�T���oy\nL���	�(�����������=D%7��a��42'փ/#�����*<nzH�e��x�}���fc��\���{yXu)ς	,��I�43q������7���:m1�F$z�b������ּ�:_T���s�*0����^�w��\��я��q� ��$yg>+��T���ڳդs�Ɉ���2�����2h���J�0�N��t�6��T�����tk�,�A
����d�}x�����^��s����.��J--mS�����ݮ�+?֍�gC^�h�R����ی5�V?F���KuV��y�Ȫ��+�:m��si�a˵��f���$&��@)Z�ۯD�AHZ!YT�1 �#��,�{��q)-��~O,�^�w��������8npS�"��h�\�T�w�l�}�M��}O׬��{9R�a)F_F�	��
���`?M�F�z4��^�Y��ֿ1=Zax�<{P5Z���foQ�SMs!e
�}P�I�b-Q�[>�\���z�U�=��h+����gx�GEA�j�����Y����y��a;7ІjvK�{�2�0{7,��-Q)xq����NJ/~���spXS�2:L���C\ؘ�jӲ(�ma��2f�����M����D�,3�T�B�݋	���'hE
�rb�޵5�Aߩ�.�P��R���(��P\�0��Ϗ��ֆ��ļ6z�GJ$E&+X�p��Ht�#Ƅү�]�A��N�ɮ�+�ճ6%��YW5}Ȓ���{�l�܎�Щu����$�X%e�Mp<�?