

#REVISION: Rev: 6
X1 1 2 V1  PMOS  
X2 V1 B 1  PMOS  
X3 2 A V1  PMOS  
X4 3 B V1  PMOS  
X5 Vo 4 V1  PMOS  
X6 4 A 1  PMOS  
X7 1 3 4  PMOS  
X8 2 A 0  NMOS  
X9 3 B 0  NMOS  
X10 4 2 5  NMOS  
X11 5 3 0  NMOS  
X12 6 A 4  NMOS  
X13 0 3 6  NMOS  
X14 Vo 4 0  NMOS  
C1 Vo 0  1n  

.END
