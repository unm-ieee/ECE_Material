*ECE322L Audio Amp - 04032013

Vcc 1 0 DC 5
V1 5 0 AC 0.01 0

C1 3 4 1.0uF

R1 2 4 400k
R2 2 5 4.8k
R3 2 8 ????
R4 2 10 77.7k
R5 2 11 ????
R6 1 3 10.0k
R7 4 0 100.0K
R8 2 7 ????
R9 6 0 5.5k
R10 7 0 ????
R11 10 0 2.2M
R12 12 0 1846
R13 12 0 8
R14 9 0 ????

*Qxxx C B E NPN
Q1 5 4 6 NPN
Q2 8 7 9 NPN
Q3 1 10 12 NPN

.MODEL NPN NPN(BF=146 IS=34.401E-15)

.OP
