XlxV64EB    2876     ab0Dl��24�wvi�������ŉ��Ӕ��b?��,��^T��'�PI����Ɉ��'�S��	�a��]��ο�+]�L�d�;l˪����W����Y�S�~�"Ci����I?����'�� �/�����HŨ����r�B���de����1,=s��_���rL���:(��o�Z_����~<Ý��X�!�R��X����)���Msu���V���B�H�k�JT�`8x��e������R#'�`V����+��������*�g�MO+x�J�o�F�`�E1��Vb�k�ݢ���=�}Y���M3��J	�Q�CǸ@�%4��d�VYDSk���7?�ǽ&�G�{S�������ER�M�
8-$V���r�ʎ��-������D���Ӡ}y�GS���\
ԣ���Ec^jΈ@y�o�,�~t/8�+������
{�7����ޣ��m�e��v�(�J���Q�w�i�|u��8�H�;N����g�Yl�^��[���GKH��S�ʷ�i���d���h�K%��췘&���%1:Z�f`�s���PA�=	�!�	���ؕW��G�b:}�a�w�M�L�:�L��<��m%����qs���
쨻S�mٕ���z��lT��}�Ƴg�}����*�������!�M�^��:#�?����;�
|����x *� u����*�'�U���s؄o\�j?:� C�Z(�h��/�ytG�f+�恌r_?�[;���1ɡ��dq���Q�~5�<�G����}�w�0C����V匏[��F�_�/�YB�cf�v �o~�G�zM���Q�+��5��!����	.QC+�oU�v�M-���T�C\��(���0U�.3���>&�!y�&:��A�%e����1.���pl��� ���t��d솰��|OT>�K�l^��@8�F5��[?J���ȓ�K�6��
Ͼ���T.3�	޽�lGho��,���N@p�,T�S�ܹ�[�oyT��H�ȷv��B�"��I�]b_ LzA۱��e~#�m?�DTl�\�XXn³������`����e���W�vr��Vħ�)�ɱ�������
��p�L����k���g�]�b��~�����]�/��kR��C��GRc��#K����N[�ʿ\�G�^V�p��V�!����8o_���G[k:�\�$�4�A[
u��K��Jw���d�	��MBf*x4P9>c� BsS2���R�N:bRt(5t��S ��;&Y���﻿��)�̶-�E3`�aMh�G��5�+Y�ˏ������m��J7���ǋV�p�X�����g]���pf{X 5�)��[*���n9���ZE`�䊙��ʰ�
�)�<C����B�E���Ɲ0'��p�����W��.@�]7��A�O���y�O��a%����/�:Oo,3}�%n��i��\�A��V�tb����gM(���Dm�^|� Q>5���H-*�Y��h��VG���'T��)���EKO�s�渕->��ҟ�!�`�<���hk=�Y1t硖:&ǝ�V�k����Ng@�Q�k��/�/]�V���&�X�e_)��`��+2C��!�<�{�Q���/F0�#��6(�x��ƴ���K�?^���y�fla�C:�9�w ��=�ۨ��>�TeK��<K�v����N)��(��֝o3u�-k�ΐ�U���U�������Q7tԾK�l��7���P���F�-٤�=6���C8|���h ��<��E��竌=9  2ŭv���%��hb�- jm��ҜDj꒨�[��x�T��x=������k蒜��H�h�B�?f��Fg�/ҎFjzm�^����A8/��������1k���u��uT���L̉���@��S���ut�[Y�D�y<!�1����h9����p��@��αL�M?[�z7����^%Pm�D�]�#4����V�*���o�N�hP��/�MovS�n�o�����#����t���FG˽	R��x>B���0���L�^jj!��l[|�n�J���L1ͩ���Ȳ�_3�(����d��B����sZ!�v����R�g�{ڈuCM����?��(K���eV���՞��#O���h�5�}����4W��e~KSi�=ݶm�&��P�Φ�+��ޓ|�������L<�`{� N�������h9�vx��x�����
�4�U##�!{UH�)��U� E�#�IZ�x��s�i�����.HY��CF2�����tt1G#��RC�
%�m���}ݟ͝"Dg5���.;�Gpƽ1�|�l��-���0���N��oG�9o��@a�A'݆b�p�=�Sl!�nK������B�I�/b>n��I�|i��6|l|�mpcf�����F&]�gڟ���������q`!��$���\��������RQ)9�ENe�'AB�~�_�@��E&����j$���gkݗ���<��bd/������ឩ ��j-�Q��;H ^��\�~��n���[T{q8�cA�='ܔ�3aǠ]�=Y������=rЌ��AZ	#�"D*��
T'^(h����Y7�.�,LS��1a�d̚�*�F�8m��ڕ��o��~M�CD8_P�Vi�$j��FH��v�`��|z@��VE2��3�O�6e@-$�a��

<p�(夜��`���R\��%EqH�g�t&� ����m�E ʀMt�u�d�����