*ECE322L Lab 4

R1 1 2 50.9k
R2 0 1 12.62K
RC 2 3 2.2K
RE 4 0 434
VDD 2 0 10V
Q1 3 1 4 NPN

.MODEL NPN NPN(BF=140 CJC=20pf CJE=20pf)

