* Circuit Extracted by Tanner Research's L-Edit V7.12 / Extract V4.00 ;
* TDB File:  C:\Users\Tony\Desktop\321_Project\RunFrom\spread3, Cell:  Cell0
* Extract Definition File:  C:\Users\Tony\Desktop\321_Project\RunFrom\template.ext
* Extract Date and Time:  12/02/2012 - 18:44

.include 2um_CMOS.modlib


* NODE NAME ALIASES
*       4 = I1 (216.999,-87.499)


M1 3 7 5 1 cmosp L=2u W=5u AD=82.5p PD=53u AS=40p PS=26u 
* M1 DRAIN GATE SOURCE BULK (173.5 -82.5 175.5 -77.5) 
M2 3 6 4 1 cmosp L=2u W=5u AD=82.5p PD=53u AS=40p PS=26u 
* M2 DRAIN GATE SOURCE BULK (200.5 -82.5 202.5 -77.5) 
M3 6 7 1 1 cmosp L=2u W=5u AD=27.5p PD=21u AS=40p PS=26u 
* M3 DRAIN GATE SOURCE BULK (147.5 -82.5 149.5 -77.5) 
M4 3 7 4 2 cmosn L=2u W=5u AD=62.5p PD=45u AS=60p PS=34u 
* M4 DRAIN GATE SOURCE BULK (204.5 -118 206.5 -113) 
M5 3 8 5 2 cmosn L=2u W=5u AD=62.5p PD=45u AS=42.5p PS=27u 
* M5 DRAIN GATE SOURCE BULK (174 -118 176 -113) 
M6 6 7 2 2 cmosn L=2u W=5u AD=27.5p PD=21u AS=40p PS=26u 
* M6 DRAIN GATE SOURCE BULK (147.5 -118 149.5 -113) 

* Total Nodes: 8
* Total Elements: 6
* Extract Elapsed Time: 0 seconds
.END
