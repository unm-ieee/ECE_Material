XlxV64EB    1f28     980��D`J�|��y������lj���\цهj��ns4�n;�MgV���\ׇ�w��;���나<�4R�r�*��x��fR�ܜ�8�>�&m̤�-CJr�R�
��Od��L�-rh'�먉J�*�V���DN�ÜW�8'	���H�F�ӧ����a�O��R�C���r���97I��#0��� ����yJ-J�g�3�і�������hn�\� p���9��S�L ��i�VL��l*��ꆫ��H�j������P 0�_R)ҕg�"�5a�4G=�D[CH�����:���,�G��tH�����v{���yC�؀S��+�����k�|[F�Q����8�Ձ�m��tF*Ց���l^W�7�GFQ^A�A���"����.yFs�_���hR_����/�J��ﴊu���q/	v��g����G�����DJ]QKqcq\�>���y��R�BX�aR��2�v���4"m�sm���BӀ�ٞMIo�N\[�>�#<M������"*�ݔ��o̩W�ڴ� �,�w6���9J�r������An�*�7�f��������֙�	��+��^F��ǌ���-DO��pJ,�`�/q*�}_��;�4}�����G�.XҤ��	Is&�ɇ���~��D�k����i��A�e)�Rb}��k�M�K�bg��.�>>{��Tc��tf:p
ފ���l>�ƾ��M�`�gY.:ɾ����YV4P�\�����`M���ocw��k��>��^���]/�Z=�RG__�j��)RI����N`W*H�Jy^YrlI����<Ԁd&F�]�	n�]���(����	�P���*�����v>��ʫ�o�JW
���D��o��k�$ƅP�X�����`�����0.����Z}����-�󋦛���C�zz�.�;�5��rK`�����[�$��4��ڽ%a����5`B"+�=9�	���\r�e^���0zs`mE�rj�m>V^墛�VU�jk�?�a]��rO4$��޹[��wU�s,v]a�����r�?���ϵ\�������*k��O]r� �9���
��O���$Lc���bA����m��S��]����W�	5�� �U1�Vb2��,\�r�!�${��t�Z	�[J ^��Dfخ������L|�)��+s[2�p�XU<����k���d@�s�`�Y���/��@B7=��?���d���JIoZ��E����[�5d���56���j�Uhj��r�u� ������fb��I�)�[#-Zd�y�M�=Gd��[�}�fpS������P?9�ؓ0�oͨ�=O�	i2ƪ�5����}�ӚU�کɆG��r'�TC��r���� ��pK����lEe⍚��]�*@VXW�EU��\�J�m&�1q����}��������~���=]�҄j���΀>����c�k6~�UE��$F��@j�;�+�����_<՜D'�C�
�g�lE��v5�V��9��
"_���>j> �~�dLȻ�k`r�	Z��f�6�V�5[кqS��]	q��
<�j󜊣Do�Պ�\9����F:���	�i,Ż�5R1M@�^�/�P&Ȅ�K�+\�Y;tJjP��ӎ�δώUX��D��� ��K1��`�7T�x!�W�#i�p�Ԑ���d��!�=�֋�FS�8 ?��$6[�ӂ`���K(yH�q>ޖI1���)ED+���R��km��s�En�'K�Z�]���mqG8?�6�2?�'i�0��d/��,�e��3�Gs�Z<���L�,�b1I"�7z�Ӑ����AuW�,TC!�އ��n�|� �J�qM8���^�4B����Hd6���c��0�)��ǎ�8�qU��}��򑹻��z���f(_NH#��~*`Y�sy�2q�Y���+%Ӱ�Վ�ѷ`8�\��lg�~�z�dT� ��&l6��J�0!{�q�-?9�Q�����஥��'7x��&���&�C��dt�J忝N�Gગ9�Y���:@W�f6�T\׮��3X��" 7+Ȝ���tK��������'�k�Q�;k����^�C��ɣ�5��H_����lf�g�vҍ��µ���R��I�B�A���F/�Vq|��jA�c�rN4o�̓��i��� �)����Q)�N��?)��;���	��S6[
_(F���?��_�h2.<~w��a�i�E=�i!���u)��X�y��щ�Fd��]�o�C���X���Aw�����K�-�����y�L�ȣ%�vP ��4X�5�=�tm�re.���}�XYل&����rs6@�����]����V�-��#RN���2��+dѪ�i��N@,����C���%9�&�쵖*������a�B�n�N@�e��T�?
��