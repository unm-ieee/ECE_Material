XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����/pខN�^H<
|F�\�
�&�0�;���+Qkp��~��l�/O���ʈ����QҔc��f��-.�2��RՙjӸ�����Aj8�O��D����WBl�KA����N�p�:�v) 8ն�������?H.��'��#����;����^�| H�Fl�ʖ�崌aA��/!G�f���Q�D´ �}PP�����~5#���El��0���4��x0�U�3��0�gS5߻je#�~�m#ڡl��/?=J����Š��e�AB��ڿ"�(6��OjC|u(�,%�G����3k�t��ϫ�-���W��������W�G�w�IȾ$�8:!��=9�-62�h��"���uz.p8���>��H}�L�X���`��bx��()��n�dex=��s�d�������2[�a�ʥӭ��(no<��Rx��@�Xz,����9	[Hr�H:M�^����Qd���Q���s98��^1�P���J鐒/���y1�r]�1��ޱ%koz~W�7��}�����f�}�Xʽ}�L&��|��	$J�JH�ܒF�J��oO�Q/�~���ZyNɲ�t��߫���Wv4Hh kו1�:���ƿx�_^�'�[����ؤ|����sPa<�J�\bj�t��X�S�9ԩ˺��{���9��V�`=2;t�n�p�]����;�?�z��8Ӑ&HS��s�'Y귬;,Nȹ;�V�5�ߛo5��0�������^d����y���>j��	�XlxVHYEB     400     1e0Reb����
����z� 6����R3�(�x*$r}0TA�T����h\��<~�f�쩓�P?�}�u\��/c�^OU4�?�Ѥ�+׮AI>���TPSB�kA���G-��|��mС咏*h�w��(5�1HE��@��s���/���I^g�
�gu�ݼ5�]���T�Pd �hA)>�_������&�=�9���c�J̿��.d��H���9`�G/:�i�ε�%8�'�D������'��=� �a����D�L;@>���r��$�2`m���c28Ab��|s���T�A%�v����O6|�)��s�p����q��_��"[Z����["h������î��;T�;��0dZ��4��z��m"Q��bSb�C��øTQᓩp켘�v!���a���#2G���+�%�ޮL�u�����hJ%�št� 
�o^/s�I֐��ƥF%��b�ͬ2�������XlxVHYEB     400     270_����W��{�`<n-H27�Q��Cv`daO��ҮK^�������W�Bc�F����f~�<Y��U�|6B<�[z
p�_P�w���>ú�v�f\>W�kզ2��ͷm��l}m�Ϡ�u���m?�H�kSݦ$e�2���ua�o{~�;#�M��uA����c��5%�S����ݓ@ ��z>�5<�22Bِ����<؄ڔ�NA+y���:�Ń�l��Ao��\_ê?jp�RMʴ��P��T��k6v������K;.>3�Ji�ݐPq �Y�1��$�y�u�	;ŐSF���������������
��/����n���8JϾ�u���̸@�a��rU�-������U�+��C6q9��\pL�ʳsŢz��=(��6}�	X�`�j�D�$�;?)�.L��i�lL3)�&o#�M��;~�)Ƒ�R�����&਱t��|㞛]Q.s��,W����N�ÂV�]�A2US@0�R���w�x3��%ܐ�"�����=ذM����L� ,��덚yiC��
�l�
�
S�&�U�3�[u����#��;��4��ot^�O����E(�Q�c���)ڻo�|:�%٫XlxVHYEB     400     210b����[�x�S���z�S�vc�a'"��vM_�6kq�尒����ݿ�&��~�Xw����:����\C�+~D／ �zf��n���9o�,�V�DA|�?%�Qгș*�dł[7����_~���5�b[��9�����\���-6K���N�:������:�`��}�;�t�σw��� �gĎ\`�ܟ�JC;���[�ŕ��8Ą�@�����|�M뿜���M>Y�Q �$7.������*cPV4�;'`�Pi5r�pZρ��x��__�^q�����<@Z��J�(b�>�:�p̖�tu�]��L���}�#���2�o$�����zǚ����Uk�֢'/��R7��q�$ͮ��^�H�U>f�p������2rRs��T���X�W/ь�P���4Z��ixL�vHd����Ë�E�!��c���(1Z��y��2T�TV�O���Xa���|q��'GQw��9q�*����T�J�5�#��~��8e%�=��V�D�n!�p���1��j�B6�XlxVHYEB     400     1b0�'XB���>�v�6!�R6�<�+<�iN�jx�+����>u�u�R��� 19�e`}��T�K��D�|�	�Kt����R�٣���i�!�{E.7Kd(���d�O���M$U�φw_��SR�v�6_:l��Yj�[�|���d+�z��h��>`,ȡBv)ˊk-�1�E*d8�gi�c�D
�a�����NFS��o���R2�!1�Gi<Tt��l�a)���1����5`I�N�f����8&�0)�/���-�@��$!-��C�&0�����Wd�w���M���`�7�J�>L��|e%��˘ʯ�p�������oH����Rl�	��>�	��H��U?㬱^a�2�k�7_��=r2�V���H�GR�5��=f`H����2�f�0�I��t)
�~O��Α� ��W��a)���t�XlxVHYEB     400     150��l
j=K�΂��o�j�5L$��Ph���l�3��ÿk2s�'�?��)��:6g���un���̢�H�N�3������v�Ň��7���W?�����#rM�ߩv�7�&�	�nc>��'�����܍ӥ�z4�����I?�-?X���3��T�����`U���,x��B�t�'HR�c���g��uq� �uW/[�����ȤP�e^����pe���G����ܻ�m���7����}�� �`����5<�Wx3_��9��/��2�4����N��[�7��@��h]��Tu���L��1�j��:���N}�����.�k���2'���XlxVHYEB     400     1b0ޢ�Lʢ�	'1�2+��t\�!��ѹ@8��N�Z��hgh�ҽ��0��%��כ.!?D���M������K]���h�P{$^t��,)�Lu�ca���[p�ʔeA�f%�0�RCVV�����r0Vj��dKƨS=�k��tX���;X<}*>�P�`�Eq�"f#�Ff`�X�=�$� �xל/�cwQD���7-D���C�����$8@0	��2�g[����D������Z:N�A��h���<܄i��{��n�-���V�|��ݐ��(�QȮ�	]/`W�f�T[WU#d�-��H�)�naY܊��)1:��OUn��@֐x/�e2��=��_���W��盛���$�hM��1�䌨���9��)��62�� ���ڑ���F#���v�
���b�QKyN�^��7x��F��n�U�XlxVHYEB     400     160nǌ���;�#V����\Z	%��@�F���u���ݟ3^PD��}w�!�ф3 ��р��ܐ9p��HR/��(7P��[����o,��H_��xv��v�lADG"�޻�.\��gz��XWSL��m�d��g`�Kq��'?T ��f�q�${0S��MNo���)s���ڲ8(�s����o�>X��{+�x
�s#z5�nל���o�:�sjmYғ�2�0�H{�ϵ�˶>?g6Ѡ<iSMF��M�вj��m:{��|![c��1�z�.|�N�f<�Y�B-��Ƙ�p�9@��I��(���ԗ;m�5���5P���	��U��X�I2�p�2XlxVHYEB     400     130w��2#��j-�7�K�U'n��w�Z�c*�[���(oyls�'�/l�G��C)��4��'�c���Q�WH��]oa�Չ~��vu���33�q�-n� �*��'�xv	f ���$1+d,h�+O�w&�w�i��K`���Y�R�c�����.��"��+;�� �`}��$�:^��=���Q����m��ו�hC�\�=겪��G�9!���eq2��ƛ���V��D��b,����"%�X7W�p�%'�P��z�{ӿW���v����"/w�R��*�دf�15o�XlxVHYEB     400     170�g
m����͊����2�;�+!����"kq7��0Iv�X(� �R��A�s0���t:�1�8wwp����,A�к���ꁣ�\@J�q}{7�ͬ;bq뤜2B:�g���p+Ԋ}B�/��]��>9̷���|UG��ܪ���q6X狒���4�dlb޳ ��D����7�O"v�`�H�vK���<�B��� R����r��am�l���� �����@x���,�%���7�1�&:;>�8��T\�z1��`����EE���#Oj���>{��zn!N	�^���tb*<��H�ݹ�F,��h8fgM����I5���-�� 8mJ��.�Nw�+��JI!<T�բ�pJU=	�XlxVHYEB     400     130�W�M�m��+-].�n��aj;ڋAo9u��|��2�Y &��}�3ugܘJ}C	� ����LRH��р	U'�H��rr���C��iS�ק�h�t�s:ҡډ^c/ړ���q|���q[�%���R�X��� �����/�b ��i�Z�~t�&��vV}��OF^aH3|b�oD�/��o0-"��Y#�i^�����!�����}�8�w�(7p�6UU%��&l�|�; Ae��i����u��g��*�߬>��6ke��cDU�i�\E;@��o��d���>��r�c�> �XlxVHYEB     400     130�h�4���I 7����cD4�.W��a����"4��n�����} �v�,MSJg�ڕ0r�~
;����B�LW�Z�ŀ�3�v�>�_.� q���e#L߹��=uH�2l-�QFr�^h�W���$ -�_��-�T�2<��]D�c������Ӣ�B��o	�%A�i��:k���ǯ�j6��y	`]���_��X1�2��l���N�V�:��TO����>X��?Gv���xe���wzC/.�� ����uo�E��ڂ����=�����JX���߭ٳcw!��<��d�D3Q�A�IXlxVHYEB     400     120�h�4���I 7����c�Ɇ�Ha�#��[�Y (�i>m�k���W��h�������[ίE��0�*w��nI��*syH`�oh�IyK;H8���
�bdĺb�d��q�U��cm�ˡ)}sf�>��a�@���v>�M���d��� K�-�w��ƫ^��\}�%���a����a�MP�t�����i��Y��A/ּpGZ��h����'j�ڽI1��!��a�ܣ+�~���q����m�Qx�6��m��������S�w�����?'U٪��c��#I��2Z�̠�XlxVHYEB     400     120�h�4���I 7����c���I$I�F��izq���:[�D5В��A��y����h�Z���G� FZ-�\��%7���+}��lD�ƌR(�ѫF֝��2�ƽ{���`���l��5�Bp�`G���Ji+��탑�3��-�}H��4UA��%��Tƹ���GqT���r	���9��9M���!e'iV-����#x%%Dd�ms�c'`�H���1-rkؑk�ѧ��!��i�{��N�����7f+\y���ӹOj�W|6���ܢ!�hv���F��XlxVHYEB     400     130�h�4���I 7����c�Q�"ޏ�Ǘɮ���Q!�Gkɘ�3��i���GZQ��fYR4��e��dnz/G�	�c��_�X��[���G�)�z��!8Tx�����i�q�������N���Զ����#��0	)�fh��Qԣ�r�[\>�<�|�ިp� ��y&&��?0_I+]W1U�;(8K�I������u����Z$]hS�~^ᎏp|�N3�x?�p��m����#8��/	́]3�k��3Ο��
}N��K��%�4U�;��	=�� �#�7%G���<<�;&g��N�'�H�XI�XlxVHYEB     400     120��g)���?o�����T��B�0[*DB T9�"�T��W)�G
0'�P{`([��jzJj`I�?���.������hEY���M�q2dR��-�Ʀː�.��@}pq4��:l�hp�*E���ʶ<�e��s�9�<ޟ��X�������Fw�fѪ�ۯ#_��)�Q�<H@�	/���|Ge<�S]@
�e퉿|,�IyH�#�&�)�r૝{h9�>���"������)9�l����9
bI���оGڇdw�����'�yh�dQw��-i}Ť阍'ܓ<ܼXlxVHYEB     400     190��3�n�V��t�Ξ�䎀�͏γ��\W��C �˙�~O�Iv �1�W����vD�w�+!b����P��~F��/��y{
sO=5L~�b_�[��x9G�@�kj�,����5j�w�ƞ���|�O�7+�W��;箍�������vr����(,�I�mj�M�(&+T>�����p��kk>e/,+�S���z�	Wl� :Xt����A�A�%d����bI�S+���D�7���	�H|YE��]6=�̫|.�Z[���3�'�>h) ]r����
�.2���\x�k*>��+�����n�3;�:�������x�7��o�LɅ��3M�x�q�K��@\� �P����yӡ��9ٳ��X^�Y6·4��c�.�Aȃ2vD�'xM*��XlxVHYEB     400     130ic�<[��̒q�|
oqS���:d+p�ݮ���]�#�5ҏd"gB/֠'J'���sn۝��[��2S/���ld�R�_�iֽ8���X�]ݜ]��=���u`h��(�m%jy
�s ������t՚��+jl��6�=�
@Bi����K�_�"�)��QC���C+�����7 w��>*srIa��JJ�'�!,tn,(��[q��/����yG���TD����x59C�����A��؆�o��q�_,���v l	�e�PJ�Ǐ⦧��T�iTg� Hڄ1�t���y�/XlxVHYEB     400      e0�'��q�U��K��P5K2f����#<�Q`l�Kj�X���P1>�Z�d<�����y��G�a�{������9��I^�WK�L�yF�O�g��WĂX�^�O*&�c*��CS?��~Z��&`oG+LG]���+�r\@A�\@2l>�7���N�~<�*�H6�l���T�qFv32���|��!�,�Z�:�I#�/���<t5�B|+�4�Y�Ԯ����[�;q�XlxVHYEB     400      f0n�9Lp�3�S�.�np��X�=[��T'��e�k!u7�\� 3��T%$���z=q��&�Hlv�Ah�>��1��g�2H�Kp�H`}q: ��W����.E{�{|�ډ-�+(��{��(����P{���]7q/�%��&:��ۮ���h��jC[���c��!l��3��	��nჵ���Ĉ'6�ȃ�R�y����]ޕ&�:w]��Y�yQ5��T�,�_�;��:]N7�ʚ�x���XlxVHYEB     400      f0<=n���l32����K�[$4b�h<?ě��!�ڡ�0��~L��u���Ϸ�;뿨�=��Nrr\��`|��U�s�|�z��F���C@i�hش�cL�Ia.��)����$�	A���������*cƗS��vC�65c�����q�o"���r���w��7�n�\�9G�T���u�������7����W�\�K�iK��J�ͫ:'�W��S�d�XG5�8\ �9���h<zXlxVHYEB     400     140'8����9׳,�~�~�� �p�:H��(�Mu�Z���U�'�I�0����}D�}�?'%QYF,����?O��`�Y\(?&X�������Y�0��)ܓy���T;k�L~�*�5h	�\����?{R��ѹmɻn `P��1���Q�������-���C�%��I�������bTD��mX�=���k�x�ᦄ~��Y^�b���]�*W,a��"~"�"�8k��D�~����h���W��H?6S���|���ʜua��
�>SI�ݬ��3�y��։J�+�c��U�]8�?�����~���kMO_�XlxVHYEB     400     180����3!�tt�E�R%2Z���o��B	����BO����ȵ�r@v�ئ ��w��7[���n3��j��)��X�Vo�y�}1j�3b�g�+g��:HD���p��� 0W�j~o���ϼ�)]�� *"i�;[t�x�W���I-HE%�7��qѱ t���(]�Ğw{oV�$��,
�D\{���ͯHA�7�>q�F!��֮�ylw���#�=��ﮆ���.��^��H
9��@�9a@M��F"��;���'!k�T}r��D�,ǂ�����+�LCR����EgD^Wd���`��1)$��;���XJ�s/�ǒ�S�rjsE��5z�Q)σ�p�D`���.{|�����b��e�XlxVHYEB     400     160�薘�N^�;�p�N�d�v��\����`�����,ۿ�7UM�o�x��S-J:�WV�/�������-0�&CU>���<�V�*����LӦy���B�g��J4�5�yC«�oKAF�tsmD��N�uL�m
\\�`��b~��/~��7�Xn�0ϬV�-���`��[tݸ��������~�@{�1=���j���ϰ��K{r�D��
��E�V
``��{2�/s������35:ȅ��"L�1,0�V�܆��`[��`6!>��?Su'����o��eR�Q�5�TM�����p�M��(�(/��F��3#WE�I���	g�pi���>XlxVHYEB     400     150j?��(��_,_4K<�[.a��&4ʀ�D����6ϞY.�a�4ZV<��
�K���"�=�]��G��0O��}��X�~�c���B���4��^�C�)ԙ��Q8[YNx���Ɵ�
_�ꊱ6��?U3�A�p�Oύ�3rzݫ#X�-)�9�V��з�=RQG�2�s���^W#!��ʹ��t�ϋ��K�R�\�2-��/��@Ѭ��Q!���3�b��(�;����JQ���'���C��{�P���Q��L��V�}~.�W������j4}�֯Be׹�G��wtz��l�n�E�R�P�`yD&"����I��EXlxVHYEB     400      b0%\�5�� �_��lA-׼x�m��K�̖��H ��AӹÅ����ވ��T[��B���Q�&�w؎��(+4�΀��@?v�Q�핹�[
�n@~b��x�l"t�u���\,����E�=�x��4BVOGH��5_v��c5�t��n}�0�e,���,��X���XlxVHYEB     400     150�ij�z��j��bYo���wQ�0�*���.����P��L��,��r����B�05em"Wğ�Oà�RXk�i96Sel'vЌ�M�rI5?R<���-�\������%}�Y4��@W~�ᢝ��4s<D�?X���b.�-:H�4�o/��W�M9�]�.�ږ��|������0T$T�~��6�M��#5��!���r,�#t4%$�cm�Q�r;����#*�Ke�5l]f�L�C����tx�T��(�����;=5��+�	���oJ$y�q�V��k6��[��?�c�&N��1
m���n���v����]�Tzq�q��� D�XlxVHYEB     400     160�@�����.����a���L�����k�����S� ��J���X�@���*u�l�L)�^�U_*KĈ�a�������)�O�S;럔Ѐ2*:rj�jlN���A(z��xΈ(YA�d�
f�Pn�p�%K���>D85w<@��C�҃�􀧸;���l����ݘtX�H}�.�v1{�����B�,�����<�H��*O�����f�+��%�N�:�&Q�(���H���]�y�ci��|��Y�)j&�b�8K-1���������o��Q�NS����o �2�:g-����s��L���yס�Y}��f�]Iiz�uY@R��=���/��JP5�]�#�z�����G���@�MXlxVHYEB     400     170�	CEOv(��
��by��_�d�E�fy�+q��@�K�^��P�/���`r�Ӗ�#C�lS��+�K�p��3�L�F;��R�"�)B��\�d�ӕ*�P��Қ�Unڪg�/�R��hs�����$��İ߾GEU<�q�G/�9�������``ڱ�ro_��x�I�������q^N�o�wM���_��Ԑ4�l
��ᶪ��Jn���%�ʭ$ �0Mؐ�7 
"25�F�x��s�QD7�XV����XNhP~������_P���Z��o;È�1����Y��$�FO��i��H8�L˒�����Y ̗���	�F>��>�8��H�F�Y�w$k)/cL�XҰ����tJY��IbXlxVHYEB     400     150wc b�A���� ���[J&�0A�YW�;�M�j0�6_Eɲ8�'��Ӏ���Cױs�qr�ƚ�x�;�$T����F���tR���A>};������mۦ/����'
��<AlflӠ[Q9]�a/t��QBͦ��Aq�Zl��E1����?K�+o�F3��Cu+x���{�&���d�.�S�,i[�Ȱ�'�t��y)����p��$r�<{����w�X�����&=���x sBj�g*����2��!��Nӷtz���R��J��������׆㒙6��$�yw��{	������1=�� �V#�kXlxVHYEB     400      a0�3'E��i��F��/�	�,;��R���"kM�� ��ƀҩ��Qyp>F=,O������k���4J+F}��@����C�ɖ~
8�&97gW
�n�.y�	��;�x����IDhN����#���v޹�Z��!@������)���B����XlxVHYEB     400     130���>,�c�O�	YX[Τ��@���<*���<|gDuFӵ%�-���CsjY�'չ�Խ�a�$�iH�!9���!3A_?}Hm*3E�{܌U	�z̏�$f��k��W}im�2U���:���]�DEݥhGe��9��5]��.��zw�ha�Q}�����G��b�8Flc8J�`��n�g�>P�EFݥtH��Bt���h��;9�B�%�2)��=��]A#Z�) �g�l�D/q��_\��Q{;}δdY��N|gl��So2�9�|r`��_!���=���M ����P6�c�tXlxVHYEB     400     170tfzQT��M>����?f6�ɡ�!���K|<��Q��g]d�&flk�
��3�u�=�8=��<-�Ky�4�n�E��5�0�|a�Ѧ�ڕ⌭��l5�f_�Lx��e�ӂ�n��	��ܮI�� S�E��uL��S6��UO
��Bc�����0�W��7�R��Cy,s�����{v�3*n�]ԫ{Q�g����Ǯ�wT�sE�h�����~L�R�Q�'Ģ�\��ԃ��ؖ~D����x@�F��։n}�zS�9^-Qe I�TS��Ҁ�ٻ�?x@�"�}�8KM�|�5�
�5���uv# ���f�lF5��/<�0����r��]ÿ7�a��ERl�hV^H��|qTXlxVHYEB     400     100���� Q�֫<hhEIG�V�	�Y�j�,� i����t��J�d�1Qo�:�G`'�t�5�A�2�������t��aDX�E�АG�p�b�y�\h�D=��7EZj�]B.�%��8y�i�����Լ(����L���n���])��<�^̔7�D}�g����?�"{��W�z��Z��%s��>�aJ���u�>h�w������C�_�L�Q�$�i_e�6)�t[�&�������5x�~�2��#���G��XlxVHYEB     400     110*�q#�h���o�������Ȿxv�UpPo����z�[L2 �!`?IҤ�$�_�XFo
U�HI�C�Z	SW
��FA��׆A�#txk"���W0b����/�7�`��6mbA 2�'�"o"�Z+�`���q�.���ywF�=X*�Ԇ�jؠ��>hc�h�����:��!��Lu*�[⢼	���9)
����D���6v̤��#t��Y�8{N�.�h�`URO���S�,3�ȣE�nȋ��s���zj�>�_&��$P�N�'���XlxVHYEB     400     150�D�� ������j+�I&�a�0�����^�ݼT�#O{������Z�B}=<�	0��-���_D#��E��v�V��(����F���+��?w��y=Ӂ�ϸ;cمX�P���]2�k�~����A~���$:�}����һX�_b7+�O�Y�C>~�g����0��ab2�7ݴG�!���1�r{&*�5kZȫL�L�e��ټ�B�'�1&�9����P�pK�{GÁ��\��G��B��F%�Х����4����Qo����,�j#b��G"�� ��II�_g��Qt=N\.t����*[��^�ԥ�ȩ ��*�擳��XlxVHYEB     400     140�y\�I=ї#	�q��d&�ZyA�k9+.T�8���_K�"747�(ox�\$<�����	_�����I���>�\Q_0"���贤GB8�3Ю@��s��}b��O��ʿ ���3G��}#��j�\�%�&n�)
��x����)bp1��	DI���#M���!I�c�.�R�1����B5�ĜQ�X��=T?2��|Q95�I֨�FDM�/a��<�Bt�*��s/�_��=��I�H���[��������] \PAŜ��4����{z˔��қ��L�������Z����7���`��1�� O_��=��XlxVHYEB     400     110�d����y!]���<1N�H}�t��E1%�ٚ.>��@�Ca.c�2�;����q!��
�p��:�����b=��V�>��LS!�z?���I���P̦�����}U�bսq4?��2u�VO%g_�rWӉ�Wu(9�d34X���и���B��:��־I��X5/�[�gx���TJ���&�@�z�0 ���@�d��2��ui"�ݗ�$J�zLo�]g$|��LA,} Y[��\ߙ`�pH��	?���E�;@����w���t(XlxVHYEB     400     150�tq>M|�Y=aw���-�(��ǭ�p�ȷ�KemJ�r�S
l �D�}_�
�1V������s*ȵ-�)���O�3�Jh�t�1�iO�_���|$��En݆ �Eb^7�,U�)��Z��X%f�j_�R�k�WYex�3�}_g�^$����w1��a�����yu��/��䵡�p����""��+ᳰ�jV���1�4���K�	`�;B�XZ�R�1����|���f��N�q��x~�k�i!]��v9��(`^sakq˳^�UMq�|k�G+WM*��0n=_9[27� �)���n�7�X�R���?'P��=�d
�\�L���UJ_XlxVHYEB     400     140��!�c�
]����l�,8�RD���iۿ����,����z��1�|]ʺ�/ҁ��<
^�N/�}���B"��͚
b��Q��R5�������Є�G� j��B��]�����=Z=�1��nb���g;�"��c��B��;>iH�<���h�X�L/vÑR����nZ��=�M��ُ؅��� ���K�� Q�=݋M
�w:�R��ޅ���L��~
f��')~k���H����W�V|2���u�m�D&�{-K�Uf9f9,S[�w���0�:�&f�Zv�r1�G��B9B𔧁��>K�XlxVHYEB     400     140�o����ɟ@�/�@�s�����c��}�Ԅ%m�Nl����U!Uj��ĬQ3��S��A7ïh�#�,K��|E��c邶��f�_D�#���+xP9C�c X�C�2S�TD��,!�-�80O\�4r��d��/�=�����f�T��㯏���ހf��Y_��cQЕV��7�����.�l����2�S3�l[׵?�P�ИT�]�� Hz{����9ޝeV3A:�L����6y
''(�/�8��$իP7��tw6b��q�P��P ��W�^5�G��R򤁺�a><:s�7�'�SN��u��T2�B��56��Ǔ�^�XlxVHYEB     400     190W�L t��KVV{5��ЊQ�~�˗��R�����I����0��3o�.������n�R;di�H��������{,�V|#d������0�D=	ӷ~
��p�"�a+V-A\w��,����4�TE��K�<,A�JZ���}��3���N[?t�{�����j),66����h��Ѽ!�*-%���g��ï�
}�C����w �H��V�� !v�<�־�"+���|�����/|�.L\s�D��3�o��S�U�.���z4�5�:�#	9�?�)2	��5�A�ݿ������(;�e���>3K�{��q�u��e��Ӏ<�n1��`�V��J�*�yG��Pd<��_���/��(�70���'��V��{u��r�oSD�<��̽�b�XlxVHYEB     400     1309m�Z��Ϻ=��)H�=c� ����1�	Ŏ�����SC`ӮW3#7�AaC j�	��,���G�{N⓸ң�B�{����Z:��|�d�E5D�
z�+�|/s�%k/�2��'�k�U��FX�X���s?���1����'���P�c�}�(a�S��珖�3mэ�d�d�,c*}D�7֓�S^*�<�N�!�ᓊHI9���f!4�=PE��u�\�u'8.ܲ�v Tpm*G4@r��v)�8|��ܜq��}ā�(�����S	�7�h�}	��+�v�ce��fc�Y�[�%����ޙ�XlxVHYEB     400     110�(?����N
XYyV:f�lq����*���bI���y�vY�v���������c��3m�y�"P�ih!�AE�-�.@���5���r�V��������p���%����z�D��lv���vP�?�����,�QJc[愩��U7*L�t�`u[S�q�N���I:���=c�m��B��%��e��|1���S��,bwZBCs���F����#�6���s��+]��L�p��	f|�V]���H�j��8?�&aW.���*3=�6c��XXlxVHYEB     400     110?���ɺ�㣉��8\�K�D�s��k3�SJ�]��a�<��܇�u`{r/ǒ-��7�<��ޯE��r/K�9��,�w�i <^��,"�e�oи��{"IG`+��F�<Pa��������&�_���W�#z>@�E�n7�׾o1����:�戏��h��(`$�;U�G�,�9�v��#Dbph>1�!�7�=4�;�{�� N�G�����u�k����p)&ʰL���fΔ�(�����NȲ����>�X�v0rP��C�<?lI"}XlxVHYEB     400     100TEnةf��J~�y =]�8H_�g��W�5�[��err��D>y���J�w�Xr�Cˈ�����^��tW0N>���������9���InZUq���xF�L��p�Cw�@*3)|g���U�0,z�&��	:䴤��C=�p�@$(؜1 �M�f�cD�Gלћ�|��U,7V�Z�s�e�+����,����Cc±�0���H����\�5���9ٚ^| �)o���l�)�II��⿮Y���|��pM.YXlxVHYEB     400     1101���w��F�@�#A�<�0;����nM����3z?��=�Sݣ���V��C |��[B�� �+]��`��o�_����jw�Ji�į�����7䑁���T�I`z�J�q��X���O�'[�~e��G+W`�=u�����A{�{��Zs5�Dވ"#�LȎ����`�5=���y�!f�<<\t��R�R�[����J_z��%Y��f+����w4�1s?a�T��("<����̣�/��P��ru!}�$��_V�SU��(XlxVHYEB     400     100��C\�z���;�c��q�������6;ݮ@3��b�Kڥ�%�������7������	y�h�^�Y���3wB��E���ĥd<��Θ�Ƃo9;#m���ؿ��,�P��h_���S;�<hu):<�p������ĨάvB�r�o�M�=��{:O�n*w���c=�W��������o�'��e��6
n|�a��?��{�Y�Rբ��g<�=���[�x��y�_��N�⧨��W��d�Ù!��XlxVHYEB     400     180�W'���)YѠ��C6c�-���,QZ��$A�x�:��	#�?˭��+�O�Ϙ=��	NO�@���h���btO���[%�U>����Q�Lx��h�c���6e1��Z��d<���uÐ�v�7���VQ�(K��vx-����*��08���/#P6N�*id�Բ%�:x!�C&�k�0�Jv��o��r�]�;�D�Q��E���@�O ��N�ܶ�)���߅3��m/��L�H@E�*l�Ԡ�!�w�� !/JH -bb��ΊL6��)�F������W�n��f��!~���4�q�����U
8���yS�ɡ,i�(>��hz6܊�c�3�1��2���d�|�9��4���1:�XlxVHYEB     400      c0Ve�u䇮��¥Έ�jsVC���kT>\�V}M:<��z[��JE^N�޺��}������W�����'E�S\�`��yo�Z��U"��KTS1��k�h��w�� ��KQ=r���WЬ-Q���"X~��L�]#T�52>�m��$o��_�J�G�q~)�����W%�G��� Q�kP(�>~/L�W���XlxVHYEB     400      f0[�fP�
����������1V`ȱа'��xm�C��w<]g��u������IQ|*��Hy�V��i*gX~DSr�Zu�ʎh v�1�F�F4lf@�WF]^}���P�C6������Uz����"�JWC�#�ӌtM@m���I}�/�`H�c��7[�s�Ҹ\\)��We�vԾ�����l��6iqy��<��|��B>'�(��Kxy�����Ðc��xto��|D��o7ɎT�S�XlxVHYEB     400     120��s���� d8�{�`��~�
���eai+^�v��!���+���P(B��dm}�K#�^�苶L}��ꅹ�%4��{iTQpfw���J�uxY��HȦ�t���!���Ԝ������^ŝbj���	�s|*6Ae��o=�mՈ�j3w�����=�X���e	�)	�9�'K�[$j�>5��˓7�{:�Ȇ3l`���̍&lHx�� ?`7�G��ꊹ�7�-�H�фm��,�c()P(�o�$�YF��7���
���*l#��tb�m:XlxVHYEB     3ab     140�I0nigf8Ka�@w�2�$��L����&*���fٮ����Y1�o����ov3Vj�n�Q	��³��F5 .b�TI���nhn�w�+  1�8_���/�B�/��JӮ#zVL���Dr���������F Si[�a0
�-,y��\�����nT(��h��[[�8t�m���C��'����E"�k�@�u�sq���[T�xՠ�Ⱦ,��l��z�E�.�A�{�K��0�������6я�.!>8�)�f��]�Ф�C�H�D��uܠ�R
ȵ�]��U9������h��g����:�+R�k�4�y.*�><