XlxV64EB    fa00    2700�l&j�~�8C��)�d��'#�����}��hW�h[2�M%�� ��qn�յ�Ix%�x׿1��T^p���R�uVs9KA�{z˚��j�lŤ�$�����k��BM�i$ϻ�,��`Ӄ�VD/����Xl*OGS-��1E���zdӥ&*k&$A�8VcsIj^=�v�Ҭ?�25�O�P�ZCN�G����j�� ���U��{'�_8��&~ ���:�z��}B�Q*��esk��90]8>�����Eȵ�'�1�O�}EA&�^��`p�����7�Z�V��FPjm;o-KQb�c=���2#S�@tF�+�R�y)�n;N�d�Z�KP:�t���V;�ۻ>F[��s�"�i�g��V�_n�
t�U��3~!���H:IY8�}A�f;��!-��I���x�d��N���~�E��Sƻ>�,R��d�+_�<�e��_6ȳS�vհ���������
�+X�$�|A{�lN�7BLC���Ⱥ�Z$x���6���aU�s2�O�]���u����ohp �<I��oF��N�mA�uf� F8Y�[f�x�vPE��i����a�黧�P�3K�.2X`J�۸��
 >� ܃[��� ��:A��鸣;-lh�����3Y��|I�J���sɌ�ꑱ;�}�����b.�3r�{�cyF��u����H�I���	�0�/��w�qb)�����/t��3�Cg鸷{����i�H�򊪭}6��̻����m��@�1���cLʆ0l��6�w��[��������̞֠��B�3�/��Y�́�e�YK��ΆY�q�Bq��@2�ci���a.�b���^�	�`MYj�x'�ֺN�l
S[{yu��<��鱅98�B���4Q@�c�)�P������iC����;�SD�b�+ ɔ>�w�ƚ��~8.J�����&�������7�%�Ξ��	��y��n���G9�=�m !N��I��1g�7Xj�HJ_q�J�g6���ŏ��O�v�꿛�d��69�������}(�� t����N�^"�}�i�}�̹Fj�9�Xv�9�.��g8N]�Mº��0�W�k@�^O�	`<	�� (}�&u)���1���z^��3��v���%��h��˸�(<��}��Nϰ(�i�%��x�%F�t#^D@���3���e7-Wkin9�X�{��ƨF��,�w+���M�s��G�x�8/���J�5��i@�OD�~�IU?���R!X���E�ˆp~�y����"��g�Ԁ%�\ ���k1�Ƕ���غkp��$w��;��������Ϭ]��_>m"���Eͥ���4�鋬�
Ƒ��O6�#+FQw�@�ߛ�w7�]���0{�Ïf�BpQ)P�B��2��÷�F:�����`��to�8���惷�=��2�6�`I;מTCāc��6�fh�mg���("~D���2%;p�kY��\���HTk�&k�嚛�8d�0�[���-�+���`�$��V)&�EC�1ֳ��=l�g�z$qRَrB}hH}���#j�O�|����Ws��\�g!Wz6�R�s�#1+{^�At�_C��� ^�患��غ�\(��ŷs#�p=vנ���T#&ݧ��#촠���B'lӮX��ZI���N�?�ǹh�4��wx��L*Ȫև�k���C�X��:I�<��	�7����-��lŨ&@���X�YA�m ��,��^��.���V�	yG�]7��ڀR����ytj��i�l4�n\"1��5��Vޠ�7��wI0��Š�߻�WBF�{��n=�֜c��|�P�f�\���PDn)���ݎiä㠷�3�|W�E�1�$�]��&�s��g�NY>2���L�s1�K����0���i�:������8���i�/����t�toQ�Qk��m���e�p?��:�j�k�J_���l4�_�ݤK�_t���+e\��Y�p��$ �c^4_dX���{��~Z/��yÖזw
��ޭYScKb��鄫e���'�8o��j
�M��F���Ӄ^��x-a~��g��yW�X|b�Rl�pԱ���կV�S�x��XNd� h��� �TY�z�����5&��Hb�e��r�K>��c��4����OD�.�(b�b����� ��
��Y"��HN}wy�(C^�*��(1��c}����j�=a���y�݃l���4�I���}�N�+v����� �4,�^y�E��X�(�ɩRaH�\�q�=ݠd�J�l��&��ҏ�US�s������r k9i���۱�[���������\\i�Y2��6a� ���6YJu���K,Oj~�t%t��i%�Є5&>#��<R�w�l��k+4:�/�p�"2*���MH��������/yH���։M/�y�M�Ŝ��76��nlu��G+�-���?��hF�=��fU�l���Yh*���|�eA4��i�E:��T��{Ё�.Y�M��B�k�7�<�Kފ `*5$&�;u�Ө�R(����?_��7��v<2g�&Q��C&��؟`�$"0�>DV��J����0eb;Ȁ�������O�|�RCj����a??NT�h��A��D .񖴎b�.��y�\w���������̣�w/����h)L;��I��k1f_v����m�à�6��q�T��z��|Y���Q퉰�Rw�B��s[RЅ�?�#���A�∖7��!��h�q����:��� W���c���3�O=�Y�Sr�;|���gd���PAAk�_*@��~p}.�&o��2�q�M�V��4����~�*@2	��۞�C&��ۤ�?
Q�s��7Cc��	�ma<�M�X�"�9ʏӻė��f���M���{q~GB�Rn״/k?�&+�73;�J�%���\>�pА��ԛ�
-Y����v���ۯ�ک�`l�����(���{�Oo������r%�\5��y6Ȝt�h	���6U�alկV;O.K�?:,cC�U��©���y\N���j�Q��?l�2�xPژ��NY��ɗ�ؠ���kh�1`�Ӫ�ްc�����}��4� �lPh67���w�S�N�O^?�9��O��B3����i=��e?sG�V�h�޺�E��x��� ~�YV_l�g�eŪ�ٙ�uc����\��Jn#ř��+=bSvM�����e��h�<l�>q����=h��)h��a`K�!�5���%�%���
3֏�%\h3�p9[��֚��pM:����F�U�����D~�!��Dp�ƌ-{{{-J��G����W ����e��>��b?<e�:�M6R�p� �`8�p�';	�~��^�p����_��# ���^m/=�E�3��r�����WXU&�LTqKݞ?	�U9�ߛ�𮿕��];�[>]�R�$����j����@��(��pz�m֦^w%��b��MS笔G7�%��f��Y�E��ѹ̽���%��4㪋ۧ��Q������/K�3���0h�U�	�
��V�^D؂h%�uġ~���x�d8�3�Y봄�C2�TK�S祛�.e�I�g��ڨ^ۛ��<��0sJ	�>W�fj�:�;Q�S��n�.�DLɃ��U��q:��50�U<5 �U�,��k���k�^b�0>x7O��]��k��s�GYp�]�h�_�;<���>1�4�n�+l�k&���pX�3����+����7e���5h*�ё��-���/�;`�ZP��[Ġ�
Z]�J�xA���|�k  �U"H�32%h���J�dZW#(k��1o��W��Ch�Q��O'�b��\������������(�_�Ċ��ko���U���v��d�^K�G�����᷻��Y�=���>n�7
��$�o�=Ё�[%� �Q�'`X�����H��6��ysr'֨�����(��v��x�U.AL1�5�Ռ���u��证��t��nþ͇ش!ཱི���.����7�����A@�˸��-!�7�auf���SS ���̄Ã�stbj��Ml�E8n�Ҵ��o�8�u�̙��/5<��+i�-t��Qdd�[0��t��Ϗ�h.C8lg��D/�X)�9��a�eeE&����?��@Ɔ�jR�J�VL��S�,'��� j|¶y���a�X�Z�ɿv
6}|�x]���B��@�E��!_��w*��X�fe�;�~w*d�0|-5�F�ȉ�(��1��as�Й���:�C�#�V��@% T�� A(nQ�ڀ7���y��E_k4t���V��J�~���`%#�*}���dB2�]\RЍD����č���I&����y#Px���	x��Ɋeݼ\���~xbݜ��"�
�A����ܺ��T� ��9_�ۇ6����O���i2螕en��Ԗ{��OMef�}=��Ǥ�P��� ��!��˻�.�]�}*�#�$H�w��S�䮧�ã�H	��x�(͵���9(Gyz��(���{'���\,V�����8�>��%��gq	k������%��ZD*Oj��>�T֨�I�t��9��W�&����P8��7����3$��f"-,D1���=��I�t�`���3��;e��Iq^�v��Fs�K�o6��/mg[��h��"�՘������,G	T�q��xq�Tgn�|�M����z>�k�۪L�+2�K`���@W��py�e1�����j������^��]�#��������XzIVP""5-�Ѐ�MהzD�:{!	���3�o��[�t��C߉��~	 ���Ar�)yYA^!S�C\G�7d3U*�j08<zಯ �+e瞵�zo�W�RY�<�m�_n����%K��Ov�O��-�QwsCۨ��޼ �L-ovh��I���8���L�z��?�{�t�+�:v�������om��؎�)�z�o�6��@,�F@���`p��wn-F��7��lx��s	���@��5���y�e	Uq��#� [�L--j��G��P�������8��<�z,������v<�뱙�{�!��W��5��s�|�܂����h�m�Re!2��]�plN��r��ZM���6o�����iÁМ~IV�%�rq��g}S����U��T�a1�W���"�Em�a*]#�� �A���l��c�g���T��kEG��5ë���p�Oa�A���_NȊ�@@��L`A��X~�f]tw~n�A�*k�2b9�A�6��Tp�>���&q� S��:}t�V�j3�Ԃ�
D-�C��g���Ց�a.Jɘ7���^G��W/��팊6��r������@�u�v��ٲ��m���ˤ�o�7���͋ح���D��G�ߚ�e�D �1E�)�=6��[��{p�lH�������.���=t�bw����2�\V���%���R�&&`&�q�;��l=�*No�W(!̓��B�
�m���)�ދ��\�s�{��~f��<D�I�� ̘��v�"�/����,<�c������죒�q�цo��>3�/{�^�:�x�&Q�D�ܺ��Tu�u)�Mѷ������xh���AL�mA_�,d��U��ҷ�yA 6�]��B��!L��,���!�7M�p�X����h�~G+�ɳ�G8��~@��P>w��fm7�=9�B�d�l��e��7�Qt���{A�`������@�G�-Ry�cm��0�m�+wntcDc���5.��a����Q�@���d�^�<�+�>r��yK�5��Z;����p��|���"�9��ja�"
bر�o�5�$y/lG�sճ�x� �9�	��!r��B{W<�t��^�.1�\��I��km�bh�ʭv�|,�"xII�®�Y|�YলIW�ֶin��(���r�h*�,h�9� V�����c�/@"�L&G^.	�7���#���"%�P��7��0.6�e����J�Xe����~M�4ȍC���������C�����+P:����\}1��������Ú`���єY��HY>���O�3&
�+���������w&h�-����tҝo���h�n���^/'��l���,S�ǶO5��Xk��� �0B�G��ӗf;l�n��Fu��3a;��8����਀Qf4���!>@'� ��D̈́�G�F��s�/���٠�4^g~���,�CN-^��5W;�v��Gã�S����4G���涼������Wȡ����<�Y���SQ�����ꛧ�)t?|{�@��1_#�U�
��8�3TK/z3�H�Ɗ@)L����@(��!ި�Zs��%c�t�����t ��e�����ߘ�x����q{Lv^^z�#�&�zv'��u�(]�c��)(��@�t���'�g;n����q��<�6��$����CKN����HFI�G�r��Q��tgr�-����Uv����³���dЇ#o�z�2 D��\�_2�
M�&�R-0���k�t�5ڧ�3�E��\�P��R�	�H�~䶆hi���
 �2 ��N
�߾f��&�u)�n�ֿ��i�k��!&�xm/����0F��k��m��y� u6 1Q&9R�;Uko2Gqagn�Z�4\��]�Ǖ��l�T�R���v؟o��c�vC�.	��P7���9#�B���&�#�y�Pmq߅�׆���
�6`�:�x�D��%�&2mj�� 8D�,q,���J�q^�Q������9U�G©�(��ЈG����A���2��cHCݜ��O��ܔ39�K/�����������ġ����_���X��ӛAf����B�А�9�����nԪ	|��W��ᑗ*(Rƀ��SD��-�"P}9�k����1n^/�3�m��	�
y����ؿ�Ƃ> �	m������Mfp0LY|&��h�(k�d.�,6dS٢U��(��9?.�6�	�|�c��� 8���T�z�4�r<����C�P̯H8�:���sX	h�p3szgyb7�,�P%1��m��ɇ���k�Xx̷��l��uO��|/��w�j���+�\R��&V9\�����i3��������i��I����W�Qˬǝ)*�	;�*��|��O�����.�Z�6��_rq�Js��h9��kII+.L;>PI�ԾS��z��d�X=��؋��hs���e���8+�F0H�Qs;��Ӏ����f�(N�xG�8,;-�a`�"�p��������(��Q��n��8������g����9����j�卋v��7��������im8́J���VN���Us�l`�Q��=��BLT4'ٙڴU��6AA	>�QV�ˤ��3W�������t$ f3Ģ�K�q��Y)��
�h�q�	�E�Z���ٜ�F6�/�Z���������K`ƲNB�c	��;�hr'�D���
������q�9��l�/y$��Q�:x-w	�I
U��� ��ۋ��
��~(F��d���aym�c��=Z���d4�E\�v[�<f���P+�u� ����YI5^}gn��M[�R������z�O�G��g7����W郀�~���J��FE��}�*Br6M�Q�s��@Y�O;m����惝�ı�Y����#0R��*5����>�q�1�&GmE�%���7�z����VC����[���c�$�4@�ŰkpQ����]V��&+i�����hh������7@S�V�B|�7���
{��]���t�W+݀-U����s�ɿPM�̊G��$�nWԆ���|�py���`�v�Zi;A
�I���,��b��c,�S<��2V������3VN�n���f3L��7"��E�uN���y8����Yj���U�����T;�'�Om��j(����<9����;����B,k Ya���Iο+ж���4�������$�����)?ab���ڠ�3���zh����@�ʓ�)��T%;�
wqЗ�ɞ�٧օH�B�7�ye$Ť�q��ȼ۩�e]�J�-�>�v�Z,.�L�=|R�+�Ȭ����`K�)
~���A�F�P�$���#����@+�)R���f��ΌN�o[4�sb(�|X�^��pAܽ������Xa���we��7���<=�|э���fQ�Y��S�)|�WbUμ���R��e��c���r&$=:IYm��E������������8�:�bZtj�g\l�R�8��#\�4��XEK`��>��B�G��t͎N�j�էd�u�Pw}�+��kt"~ܧ���oh�� ��%gK]r�ߠ��RM���Z��
��F�u�x��u*�N���Fl&�E��6M�$����_����5c�0�����q��.>K[tm�>�j6'��Q�J�O[����4-�Jтt� �yo���U#-u|WE�^y�!�0�[ElF�@z��`����N�:��[n,LcR٤�{�N�R9�B�M�xq��XN����Y�z!.��}3�3B��ҖAz.o��`
ɯڃ/~V�Yy��LS�X�Rػ�U>���
O
��5�t\-��'��hا���M�>�E���@L�^7vٳ*���eA���Е9�)n�>]/�wS�����x��jk�W��򙊪IS,I�n�_1����ݙ��o����٨ �VR,U�X�CV���ح����� o �A>��y�� v��25��F�9�BU�+�u��`���W���Q~`T��-W��n�_L��+��)���cV��	��C�SG�	ÒH�MZ�G(�
Q��u8%�����d�����9Ǣ�뇯���ZsF�|aY���\���˅��Ըw�Yӏkx��?n��2���!��y1���=U�Y��|�#t*s���vP���[<j�	�9r�>���ΛpG&��l�o���!��~+䂻���'��1�7;�)��;��f=�l� 2d^��n�� ����<Bst���P��#P$�naUm�Z�Iϛڿ����w���_r�5�}�,i��1��A��:V����-%V����#<� N���[���a��=�����W.j:�O�BP}�r����zO��������PF��3x�&Q&n����q��R�#l�%���(�~ANɈL$p�ҝF/jp��T�P�������T��\h�d!�a+s���h���;J���K�짚��L��G����}��*E]u�	�p��;QsO3k�sC';K���#f8X!ܝv֢�FOѱ�:D�kq�C�L�,�+Sy���Ӽ�0_�?��俖��$�&5$�_z����P�,�񞋋@Y�l���hrD�gY����!���[�{:da���H��>���x�7殟\=�������1�Z+pnH$S�t-�Bz�]�6p�x"����MO��_ꥩv��>S�^�PH�B_�'�5��R�g� �NH�'���çW5\�=��/��������o���$_ʸF�Y�_���\z�7����3�P�x,hT3޽�8�.��Z	�����.y�$�.��YH�_�ZCD�����'`�Y+��nH�ΐ�,��C^��/��m�z��t�ɐ|�#Mȑ��̽�U]���ķ�]�� � ���&"?i68i@�dq�E��я��������p{u����H�?���XQ�ۗ'
E�],wB�!���a�>��O_�'����t4wW"dɓ��C2k�8��q#q:��8Y~*�+8�=�&]E��^�P����OF�P�>�a�g�,�vW�����
.'��{����빬<�#��Y�pM��q���_rN�ZxH��M��$R��)�[���/B<*�w�?���K��T�/e8�*�Q�,����EռF\Պ�"3���_^�g��rD��c �L�����O��<XlxV64EB    9af6    16c0�x��f�\���`�(n�K_*-�0L[���=��(a>��۱l����d5��8[��(��A�����	��sr�s:��P?��i8�z�O( 	c
�_Z�һ��V�^�טM��tښ�bM�;�4e�s���m��Y�(z�����>y���Q<����z��4����X�(E�ѧ2D�ψ���"f#�ʫBK�>��fa(����T�`~�mZ��L%�l'㱳�j0^�q�/D3�D|�M
�R�7� 9l9L�'/�e� E]�<����\}����c�7v��� û�:2��I�%g.��-p����� ��<Q1�Љ�'��0�RΙ��f,��+˙u�[~x\�G��&�vH[�y�ӈ,h4 0as���E��Ք��Q���_����mF�_q;ۇb�j>���A�Ȱ�2A����\l���2�����辐9f�&ǯ��mr���a$�K�*�i�M̀���##��u3�RD���ˇ�H\�5D ��Y��j�ج�4��0^B�l�g����c����K��,~�i�EJ5�t��f�x׊{G������A��Oz����:E�A��p���M��N�o\t(E�v�ݘ���P���z���8	�ϕ�"R�Dա7�s���DX�p�*V�g-�8�T\΄z��8�'`�I��\�E~c���0�@�}�v
3RA;�W]>�֔�\(�c�_6�\��p&���@S c��9����@IY���U9[��$�d0E�+gww� >�{jZ�Y6��ǽ)~��bj(Eu
���ɇ�r����$K�v����J@F=�ƄN�:B	�u)7�mw�����ZR��UrI��/݉�x��ڔt����ķ}S�d�Er�����Tҳ�&~�����D:�qu��������i߰O��9&�zJ$�����.�<����zh�;M8KU��\bmҞ@g��r�2���;�q�q|��8�)�Od}H#����������&,62�-
@@4�ӻ������=��T]G�ÁƗy�)���+�貊�p+T��tI{����)ӵk�+a*q�k���PVc���$n讯�g�a�f�>���^�Ӿ���;wȧK��|�[��M��&���R�Ѓ��Y�{0�7e�Z�=��O� 6��ƃ.��I��A�(�f���oe��{�����~t��{�+U�p�}3�e��򲥻�ꄜ��\��G Z��E5&�:>�d҉zG�6O��$�L$���z�l�oQa9�X��28'ޡ�+��p��y�%׺QRoh���x�j�m�mz���c���`�W�陌�qE<���FLf\�-3]e1��&\T���_��[���_��\»�Ćp�p�4}e�!?f[�~��7����%Y�I�T�i�X���ă G��_��M���������t�L��+�8=E-ɲxFVɎ9�n��i(K��dB�}c���C�2̣�Ơ8��o��,cw_�`���>8Z�������4�ht������S'��&�b����������d�3�p�oM���Q�ȢF���\Kn��]?4�=��X|�S��:�����G��dh6d`���cEQ�L����ގ&�Q�y��[T����g3���������@ޞe-0��OĐ^�X��m�B���Dv���60�N��G�'aM#$�v՞"�?�I!������>j�n)��!O�H�_{�rM���Ŏ3iW�_Jw�W����-X
��_��$8��Δ�`���Bf�띊h�Jy���s%��6Ђ�Tj����X��F0�Ly�����|�o [QP������(�aN׮�cE�������c���j��gJ�&��r��^�QK��\h��i��9�1W�������Px���7����X
�i�)0��d0,�0Q���e�?ﰬ��>�@a#=FSeM �����H�7��'�����%��Ny��B^�T|o <K���D+��NS"���+zV���lO�Р��'�V�?�:�vM.��%J�Պ�,	�U����㛢]��d�`^�L�����^��mwN���DZ�M��0\�x�I����~��sAn��lӌ��%�C�6s��@�+�o�k�|��9+�(Uč}.��0�@�v��{��ɽ[��8����l�R&o%o��fbY�u:�袪8��/,"Z�sX;EV�7����q�,0[��NX��,EK���`���iM��B���肒���u''����B z�:c��%}�l2���Tr*�4*����e��$Q~�t���ɒ-ڵ�fs�T��<la�:<�r��{�IV�߭Z��(��tx�x���~�F9?�]�|�*T��گ}�ү�?5��D�N(T�0@�E	h>&ܨ����tL��(�&��m�E���ZbK�(�A��k�P� ǎ������� ~˫���f{�����c2�A��Z��Zݺ���}�4������=�ix4��d�Ѻn�Ȗr_�e�q�<�!��e��;�b�E��C%�͚Dɯ<���T���u9	:q���J䮺������7�$:X�Vk'�'O�;C��������D�'��`l#i��3���]��� �?��M��p�8=�i	=�̨�t`��:Œ3@��1�$�2�l���?�d^�Eh&�Y1���*	���ܧO�.�3۟+��CC�+f[7�Q�x��>���pvR#��=k��59�q-$\_Y�_MC�j<6��ꩬ;+t(����'����̙�wg�G�U���E6A���e�dXV�Ra+J��J��ӫ�����+` �"��o!�ڬE5���=�>ŝ�x�*� �e��)4A���%�I�q��섢\����V��IR�?I/�G��N@�����jX5��b�ч�_Խ��x�&�Vo��^e~?���A�;������͍��*0��T�PGi.��/K��GBc1��0&�iء�)�A�?��<��ܠU��f�q���X>MQhh֒@���{D>��;�K���sQ��-���ʘ/$������fP`�Gni�����cHpI����Z����J}n��c��P��s�G�"P�i�o���VJ�y�U��ľԛ ��ރ�ܮ�
/��U���\2K/_
Fw�x�<�y�L�lR�%��X`�� �a� t��YS��o<&��Nc>�baM�<cF$���#n�/w�$��dW�t"�?�5Lzӥw�/�{��q>���~�Hmp�����f7받"2���@E^�~��5>:��uv��GƉ���o��I���w8���ૠa8@� �"�DumT`�$��oD�=$��kd�,|�ՁL��_n��Uҏk�5���SR#\��-N����0��(h�KZ�I��4��9�����G)��Nߔ_}3�G�qG�:H��^��>8Z��=��?�j���[�?j/�O(�ꗴl�V� ��ۜ��qX]�AD�k�h>F_7ol=	*J$"�+3&�A��@���C���j�+�]���39���
AX�lgf�A����� �Bi8dI�a'W���U�g������l��'��k��,uLW��A<#����MRm���� 5�n�t��w���P
�ݥ~T*G����Q���nЈ�+����v 6���NA2C�7���?�BE�(��rfX��9&,�8Ċ�Ih�0&��q�j��Y!gTE�ΰu�dC�����s�؛)����#�R���D2Ԃn�m�7"�V)�đ��Ӫ&j贃����$0P��o�}����f�U<��2��p�Wu�x�~~���Y��_�ض%
��,,G�eb��TS=G?ϛǿ_F[ep��+�.F��b����B7X^Тz��[�T�5C$r�ҥ'�"��=i������^~wBv�;�@�k�=�T۲�$�Gs��k��la�xߒ��~p���LE�ze�xg�w
�,����8�|��*��GҔ��m�^B���Q��X�g����x�7�@�/���S� FK�U��T�x~Cl�'m�������\H�>X�U�艄L�}���0�ɯ<@�s����d�r������XFb-�0��<�N�r��|�J�>�g������C��3~�G�E�E�o�&�Rw&��ݤ���%�`�m���m���тDH/��	�r68-�͗���2p	@q�q0�_Wq���ǯΈ�Q��D�ы���������u����Θ�ʊ< B"�w'�HUT�i5��0I�Ђ�!�_P�I�T����#E�;_;�ħ�://f��-}�rU��ƪUD":�O���'�A��1(��5��/s/�T���܁�gԤU�n��8| �|و�6�xB�UU�BH�� e�U�5�F��fkA���f���S��%Y��/��OC6��84��8N�=l������Ú����~�`	\�;�L�4iˎ��d��H�����W��K�s��W)���ع	@N������>��L y�n�5�b��PX���(��.�G��t�c�Aݗ�8����}���Q=�m[ [�AT��(����H�����۰�1eQ��h�4̵�[N�fɺ#㖷c�2w���hHr�c�T�%��g����O� d^6����{�QJ�\�s|�^
?�֦��Zu�����>�(��A;��_�UpT .�P`��߶\҅X�m�O�`�PW�V��,�`��U�{X<H��4�q��Y�k�r@��_ﵺ����w���	� �w�6D���Ŧmso�!z�ߥz2{*ƒ�����1��(��7���P��%z�����s1�2֤i��9Z� 4����3q���&�%�,�W�+��
D��c�*����z2նtrE ���<��ZI�|�Z�X���i��0�����'� �6�a�X����}EH�A��Ϙ3�Ӈi���Q3�^��:��2�:; ��v�6���}5����� x.�k�OcS���P>�qdOq�WJ�K�`'�"���
a�t��۠�	S Ph�a���y�\��S����bd�*_?��ٰ����J�V���$NA�����P���n8a�H����5$���s��oq��p0�q<�.e�)���ŏ�D�:|
�f	G�1ג�+M�+\d�up|������xe�В��]�D:��)��e�S����C�l�Vr�� ���a$uF�^�y��uv�����4�nB=��2�u)�؀�"jY�=D�(�jy��3�]�MO3�oA�����W�>D���ǰR2V��ͯ���B�Z5���0����s4���M���!�}lN^		�B�+�X�Ӿ�ԏʜXk�����Ĕ�_+�6)#��Z��aä$x����i�Y�O��J��ٕ��f*}nh�gA����~x�y�F�,u�{+�Ѵ��)P��6�I :�0�r<�5�>t�"�P��}����%`F�@�8�Q 3��"�!��[���Kq�,c$J�c8�g� x)��r�P��HO���$;n4⩕uﱆ K�ƽ�g���v�T�	{K`2���fWzF}Z��)�3uX!�^�@�5[�`�$$P�)�d��y-���b����>I��$�B�`�:�O�Vfش��-5���m"@ @2���I�q��yf���j�c�=�Z��&C@��=��7ބ4�� ϬՃ�I#��Vٞ	`�@	#���J:�`M;��K!��+*�U��b��M��ױ�4