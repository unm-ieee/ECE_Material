XlxV64EB    116f     7a0�q�)�.��Z�ߘ��>�]f�?�vzNP��"{s�Ϭ��= 15Ӣ�Z$O��`_Q9n��Wu��_1]X�Y}�;��?����3�ԃ2�g4��F�9��B��z�7���,�1Y�[D<@n�=q����G:L�;=���~@1n�M���c����b�%�t�}�>���`�����Bq���]�9��ߜ�z9v�9N�(�c�\/yw�ְ�h���#_31���5Bs�-4�V��\Xm6";��`����k��������=���߾U?�&�Ż�t�?���~�꒼��x����<�)�cʱ���]̜�&Z�K�*�B�sd2��޵�ve9��J�X������ �^��|�t����
0�e�@�����Z�8����P�u�A��O��1�&Z�����+eǁ��zSL�z��- ^���h�"x`P˙�����~)��A�Ĳ��k"�*���̴�TP�
K���tH~61�8�
o)\�¡�?��S�Cyw����n��J#��@X���~�?�%�w�����V}ρfZ`��E<�!�.�/:
�bwԳ�����3�7ä�$�GW����T�h��� ج�J�"%����ҞSs��8%��d�+7�F~���c�6��p�efԺ(%��s姢M�y�!^"�NV2�]0��{��vU�u<9ZO�,uET��o�(����l��� �sr�2��J�$����D+ۛuϑ����Qu�@��dº��bP�ћ��\q����A�v�~�r��6Pn'���c~�����;Q?E_:�^�ȏF]	�lj��9Wg
|�	�,��5���W��POZ�64A-t��Cr�B��̤Q��'(ުUSU���^�ͣ����
���D%:�%�C!<F�4��ě�rV�A���O
�ll�� ��k�[~�W��A�HG�n0Q\�(j�H&��~F�vM6�B�f������X�]/r�D�͠CQ��IA1�R�����EdvI�p��k:���&��ꌸ�I⺿�n��]9$R�]rux�I�{�G����u.,*tV��YP�LIDel!(upl��hw}��*oKt���o���qrz1��]���%���u�GI9��W3��t�p�s
S�}.v��:��o	aݤ���ң"	gݓ�a�²�L����Z�!�����<��Y��w��̩i�E�x�O��;�5�����L@b�%�xފ����Ⳃ��J����1�������6���i�A����O3����}��Qlh��>q�$O�Y��G�i7b�0��즡���}p;���$��uR489�Ŧ����+�v���@��pN�-�	%�&�����3��>�J��C�#Ŵ�{掃���a��=�l��uk��;�;�x�cӕ~��y=̣e�	���@��z�(��|�V��M��J�]E�M�׻6�D==n�e~!�ј��z(&�F�&R0�sE�W{��~%,��� �ۡHj�("l$[�Z
jW�-����л��M8ݤ���&XMAө����=of�	1�,=�O�L����o�[`,2K��#Iя�ٓ�÷$<.Wcl�*�c�J�˨�qT�x���� ���Q��W����N���_}�����դo.�a%��/��$4]�ò�БT��?E4��Uʐ�[1/UVu�@�,6�������ؽ(�����%��ԃ/>�;�x���Y�a�j�;c�wC��CV��˒��ILN�����8�mY��ئ��M�ں�Ou�)�F��يa�A@o(| Y�O�9x�	�F��N#:[��
,�)=p,�@9oV�'d��� �p���<n*՗4C_�y�ӌG�Y��p���u�o)��E�H�`8�t{���?�ǵ�m����UD���A�A~	�w��p��g�qf��y��T��拳��А^�c��o��c�