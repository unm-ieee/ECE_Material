XlxV64EB    2245     e00ͦ��,<�k�\2V�>K��3A6�?H�+aƀ[`P�.�����U}�(����3�j��5���}?>4R���� *��;����v�*�p�ҟ|d<o���u���Aiz�ϒ��z#��oxٗ��l��N�z%Kc���E#WP�w3��>5gf��u�*q{�)�x]'ck��@���O�A�a�{@O�8z.ϵ=ۆ9I��������Zt[����� G�OV�v�ДYTGR��x�t4�ꠋ���,��&��(G�o�Ǳ� �ZSү�F���r�,�[��L7�>�H��s~��.�H��t�� �vA�a� ��{�زL��2�5��J�	Y�L
���#pп6uL���h���l��FN�-���M7�B�	9�����~X����!���Tԥ}=�����l[�*�m�DcdqG��,/�H�5����wO ;�᜴x6:�%� ���|թyӎy��2l)c��Ι֙@v�$��Ex�P��l&�\��)A^��5<Șd�� J5�O@C%����GC��ؑ;{���'��0�5��L��w���.Ϗ̬��������:#��^l��R���7bFq��A�`�8jW5=Ǜ�ϐ���K3f��t\�Q/:2�/#�&_c?J�Wc�ls�R�s�~Z!�t����e�����\N�nD��������t�޷Z�l��1��,��� /OS�Z���7"d���Qs�����R?�
}Γ����Զ�Psp����K����/��}R�M�ʨod�{6�|�D��eGAf|
�@���}��8!f���jO�Ia�&�O[d>����߶�ꝉ�A+6�onn����m�F^0�UO㵿�Kŭ+k�M(��Li���ڭ�7J"T�"8A�[��R;V`���@b5zBEE$ܵ�j�bㄾ1�/E�f0{���&=[r䐛���ձ�,�6�=��L�K���3��Z��(GA�X�f���dRNO�e턗������(�V��P�Pxv�L��r���7ш�Ю�x��U� i�FC����
�r�{`vY(��#=|gyA�H���r��_�����.l]|�ej�RB�b�މ�?�d���f��8X������!T\�;�_�*�
�i	�<x���e��Ė��"5]���2������� 3�"[Adu����e-ҢB^�����D����%E�ܧ>��*m�|�+<n�o�EV$�b�n��6A=Rx���mH�?.����ٻϣ.����Y
�v��H��B���V�K���� �JK�]�v<��"�K�v����ƀW������K�x��,2���e��+���0�G5c~��ۨ�����I��1Cx�n'M��=ذ��o�uu�8��_]��5�>�jp7�2u��K��'mtDe��<d��!��}�Lq�-&�l�^�4d���Z������j�Fa��ߒ���]Q׏Zjx}�ǁ�fOB-�0����"gJZ
r�fp�1_,.�hs���� HnT�X[ϥ�^��,-��������{��F�&�	�J?5�DR�'Yd�v������ ��`b��3��i�;ֲ�f1��;9�m��|Jv�M�
;bP��6-r!f�0�i��7:�>cm��H�(���F���;TCA�w�˱�R�Lp��Ӂ�]1;���R\� I�"-�n:��G�?�R�o3�.�#���[�gސѓJ	h��<Ɔ�����wA;D/�\b|?�ꎣ�B�,"U����o��Х���� &n%xD��W�%�hE�B�	�E��O�^�|��#}F�r�����y�Q=��fE�W!io8�U�%�@C���X����"��ʸ �	��)K����eH#�%��M]Hf3Ρ4P�/5h1[�Yh����
��D�d]]�Y-�88)��x`�������U�6����ta�$�s���u�[OIZfgx�LE<C<�7 '/ߔi�v��=��D�H,��Z�@ܐ���`:�h�a���$}��+�峎�-oy��i�^�}$O���[|n�٭g���.^�f�d�r&��n�Fh���&w�m!�����J�O��hc:x�N��3�YdD7�Ѱ��@϶g�f��B�²X���H�.���u���3l�zw��!��V���YI(�,����]"/ݧj�e���c�2kj����xW���A�%5�5-3��:]a`!�v�`�d>d�*�x�i`�ѧ�Ih�[׍|vB��0���Е��d��uF&5#��H�A��צ$<��	�p��������*���3���80���z���Xߍ�`z˥�z���	�M���f�{]?ܒeyy�J�ܤ��Uذ/,Bxw���q6Sv����և�;O��b�:��Q�Jz�i�{/�bc����?��L��<Pd����l�$	rBz*��?��^�M`ꪨ��9Go��hG_�m|Ǆ���`���
�X] ?�a�� ��Q;q?w�+�;���:��ޙ|�.F�`��uo%5=$G����S`B�"K%{)�#��o���13����S�i�$*$���U~�ܩ�����	�D9�� ���zt� 8�(��|2J�UW��
_�愓�n�g�¦S���jj<'�,`mm�Y���_"��J���=��h��H&6m���|q�H� j1��t�y�L�	tV�N乂�Ȍ��T�%��=���q{M߮�Ͻ�+��Oe�FV���+^"x���2�O}!?�1j^����Q���()K��S���s��cZ�0�X���S
�V�F���C=T[9�<��Ga�����{�nV�3����c���{��������'T]��Y*�Y�^se~e�z4k?�p��/5�t?R����>B�"��x�'�,V[�I��m��cu��ȝ�Jt���nO*�W-F��f,9�k
uŷ��v�k�g�9(��� �զ�s�{�E'z���q�޿p�4��f���ϳ���f��c#��.9�4Bl�Zm]�����k���rb�-���Z�b>	\ �n@]�Q��<��/ㄚhF�ED	6����HO<��4�q�c�&ߠ@��Y����x����R}$��H춶�ٞ��naRЖE�4��}�x[�b9k\t�`T����k�����|U���av"�hbe
Wђ�\��I|:�91a�LV b�dX�g�O�����N��w<��!�G������y]�ު�{ewv�Cn�]�;f�����`d{g��ێ/]}��B�Ŕ��A�T̲FB"��ț'��h\F�{�C�'���1(_�����4����-A��1$�����71�qx�WfUa��1�}v+ET(�t��(4��d��-х�ϺF(.K`�iqh���&x�,1��9^ܑ�M��k���۰�R�~y8�U�V���WN����F/i���Ó��L��_�O:�����}:����v0#*S�#����G�a�_j��t^�ǹ��e�Ž�%�xy}�o&cA�3�=`��&*mN�j<��hf:3��%��*��C8}��Y�D�::�����s��'��p<-�/�,