*Circuit HW1, problem 1.13*

R2 N1 N2 200k

R1 N2 N5 150k

V1 N5 0  5V

Rs N5 N4 1.2k

M1 N3 N2 N4 N4 ptype l=1e-6 w=1e-6 
.model ptype pmos level=2 vto=-1 kp=250e-6

Rd N3 N1 4k

V2 0  N1 5V



.op

.end
