ECE 322L Audio Amplifier Project
* Designed by: M. Chaves, G. Iven, A. Rasoulof

#REVISION: Rev: 193

.INC ECE322L_Audio_amp.MIS
Q1 12V 13 A1  2N2222/N  
R5 A1 0  3k  
Q4 12V A5 14  2N3055/TI  
R15 14 0  18  
R16 Vout 0  8  
C4 14 Vout  1000u  
C2 A1 A2  100u  
R2 12V 13  75k  
R3 13 0  750k  
Q2 A3 A2 15  2N2222/N  
R9 15 0  100  
R8 12V A3  1.6k  
R6 12V A2  500k  
R7 A2 0  500k  
Q3 A5 A4 16  2N2222/N  
R13 16 0  68  
C3 A3 A4  100u  
R12 12V A5  1.2k  
R10 12V A4  500k  
R11 A4 0  500k  
V1 12V 0 12 
V2 0 -12V 12 
V3 17 0 AC 1   SIN 0 0.02 1k 
C1 Vin 13  47u  
R1 17 Vin  500  
C5 16 0  47p  

.INC ECE322L_Audio_amp.CMD

.END
